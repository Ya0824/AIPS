module aes_top ( reset_p, clk_48Mhz, plain_byte_in, plain_byte_valid, plain_finish, empty, cipher_byte_out, cipher_byte_valid, trig );
  input [7:0] plain_byte_in;
  output [7:0] cipher_byte_out;
  input reset_p, clk_48Mhz, plain_byte_valid, plain_finish, empty;
  output cipher_byte_valid, trig;
  wire   reset_n, init, next, ready, control_n2, control_n1, control_n21,
         control_n20, control_n19, control_n18, control_n17, control_n16,
         control_n15, control_n14, control_n13, control_n12, control_n11,
         control_n10, control_n9, control_n8, control_n7, control_n6,
         control_n5, control_n4, control_n3, control_N160, control_N150,
         control_N140, control_N130, control_N120, control_N110, control_N100,
         aes_core_n93, aes_core_n92, aes_core_n91, aes_core_n90, aes_core_n89,
         aes_core_n88, aes_core_n87, aes_core_n86, aes_core_n85, aes_core_n84,
         aes_core_n83, aes_core_n82, aes_core_n81, aes_core_n80, aes_core_n79,
         aes_core_n78, aes_core_n37, aes_core_n36, aes_core_n35, aes_core_n34,
         aes_core_n1, aes_core_n77, aes_core_n76, aes_core_n75, aes_core_n74,
         aes_core_n73, aes_core_n72, aes_core_n71, aes_core_n70, aes_core_n69,
         aes_core_n68, aes_core_n67, aes_core_n66, aes_core_n65, aes_core_n64,
         aes_core_n63, aes_core_n62, aes_core_n61, aes_core_n60, aes_core_n59,
         aes_core_n58, aes_core_n57, aes_core_n56, aes_core_n55, aes_core_n54,
         aes_core_n53, aes_core_n52, aes_core_n51, aes_core_n50, aes_core_n49,
         aes_core_n48, aes_core_n47, aes_core_n46, aes_core_n45, aes_core_n44,
         aes_core_n43, aes_core_n42, aes_core_n41, aes_core_n40, aes_core_n39,
         aes_core_n38, aes_core_n33, aes_core_n32, aes_core_n31, aes_core_n30,
         aes_core_n29, aes_core_n28, aes_core_n27, aes_core_n26, aes_core_n25,
         aes_core_n24, aes_core_n23, aes_core_n22, aes_core_n21, aes_core_n20,
         aes_core_n19, aes_core_n18, aes_core_n17, aes_core_n16, aes_core_n15,
         aes_core_n14, aes_core_n13, aes_core_n12, aes_core_n11, aes_core_n10,
         aes_core_n9, aes_core_n8, aes_core_n7, aes_core_n6, aes_core_n5,
         aes_core_n4, aes_core_n3, aes_core_n2, aes_core_key_ready,
         aes_core_enc_ready, aes_core_enc_block_n1458,
         aes_core_enc_block_n1457, aes_core_enc_block_n1456,
         aes_core_enc_block_n1455, aes_core_enc_block_n1454,
         aes_core_enc_block_n1453, aes_core_enc_block_n1452,
         aes_core_enc_block_n1451, aes_core_enc_block_n1450,
         aes_core_enc_block_n1449, aes_core_enc_block_n1448,
         aes_core_enc_block_n1447, aes_core_enc_block_n1446,
         aes_core_enc_block_n1445, aes_core_enc_block_n1444,
         aes_core_enc_block_n1443, aes_core_enc_block_n1442,
         aes_core_enc_block_n1441, aes_core_enc_block_n1440,
         aes_core_enc_block_n1439, aes_core_enc_block_n1438,
         aes_core_enc_block_n1437, aes_core_enc_block_n1436,
         aes_core_enc_block_n1435, aes_core_enc_block_n1434,
         aes_core_enc_block_n1433, aes_core_enc_block_n1432,
         aes_core_enc_block_n1431, aes_core_enc_block_n1430,
         aes_core_enc_block_n1429, aes_core_enc_block_n1428,
         aes_core_enc_block_n1427, aes_core_enc_block_n1426,
         aes_core_enc_block_n1425, aes_core_enc_block_n1424,
         aes_core_enc_block_n1423, aes_core_enc_block_n1422,
         aes_core_enc_block_n1421, aes_core_enc_block_n1420,
         aes_core_enc_block_n1419, aes_core_enc_block_n1418,
         aes_core_enc_block_n1417, aes_core_enc_block_n1416,
         aes_core_enc_block_n1415, aes_core_enc_block_n1414,
         aes_core_enc_block_n1413, aes_core_enc_block_n1412,
         aes_core_enc_block_n1411, aes_core_enc_block_n1410,
         aes_core_enc_block_n1409, aes_core_enc_block_n1408,
         aes_core_enc_block_n1407, aes_core_enc_block_n1406,
         aes_core_enc_block_n1405, aes_core_enc_block_n1404,
         aes_core_enc_block_n1403, aes_core_enc_block_n1402,
         aes_core_enc_block_n1401, aes_core_enc_block_n1400,
         aes_core_enc_block_n1399, aes_core_enc_block_n1398,
         aes_core_enc_block_n1397, aes_core_enc_block_n1396,
         aes_core_enc_block_n1395, aes_core_enc_block_n1394,
         aes_core_enc_block_n1393, aes_core_enc_block_n1392,
         aes_core_enc_block_n1391, aes_core_enc_block_n1390,
         aes_core_enc_block_n1389, aes_core_enc_block_n1388,
         aes_core_enc_block_n1387, aes_core_enc_block_n1386,
         aes_core_enc_block_n1385, aes_core_enc_block_n1384,
         aes_core_enc_block_n1383, aes_core_enc_block_n1382,
         aes_core_enc_block_n1381, aes_core_enc_block_n1380,
         aes_core_enc_block_n1379, aes_core_enc_block_n1378,
         aes_core_enc_block_n1377, aes_core_enc_block_n1376,
         aes_core_enc_block_n1375, aes_core_enc_block_n1374,
         aes_core_enc_block_n1373, aes_core_enc_block_n1372,
         aes_core_enc_block_n1371, aes_core_enc_block_n1370,
         aes_core_enc_block_n1369, aes_core_enc_block_n1368,
         aes_core_enc_block_n1367, aes_core_enc_block_n1366,
         aes_core_enc_block_n1365, aes_core_enc_block_n1364,
         aes_core_enc_block_n1363, aes_core_enc_block_n1362,
         aes_core_enc_block_n1361, aes_core_enc_block_n1360,
         aes_core_enc_block_n1359, aes_core_enc_block_n1358,
         aes_core_enc_block_n1357, aes_core_enc_block_n1356,
         aes_core_enc_block_n1355, aes_core_enc_block_n1354,
         aes_core_enc_block_n1353, aes_core_enc_block_n1352,
         aes_core_enc_block_n1351, aes_core_enc_block_n1350,
         aes_core_enc_block_n1349, aes_core_enc_block_n1348,
         aes_core_enc_block_n1347, aes_core_enc_block_n1207,
         aes_core_enc_block_n947, aes_core_enc_block_n708,
         aes_core_enc_block_n467, aes_core_enc_block_n240,
         aes_core_enc_block_n232, aes_core_enc_block_n196,
         aes_core_enc_block_n195, aes_core_enc_block_n194,
         aes_core_enc_block_n193, aes_core_enc_block_n192,
         aes_core_enc_block_n191, aes_core_enc_block_n190,
         aes_core_enc_block_n189, aes_core_enc_block_n188,
         aes_core_enc_block_n187, aes_core_enc_block_n186,
         aes_core_enc_block_n185, aes_core_enc_block_n184,
         aes_core_enc_block_n183, aes_core_enc_block_n182,
         aes_core_enc_block_n181, aes_core_enc_block_n180,
         aes_core_enc_block_n179, aes_core_enc_block_n178,
         aes_core_enc_block_n177, aes_core_enc_block_n176,
         aes_core_enc_block_n175, aes_core_enc_block_n174,
         aes_core_enc_block_n173, aes_core_enc_block_n172,
         aes_core_enc_block_n171, aes_core_enc_block_n170,
         aes_core_enc_block_n169, aes_core_enc_block_n168,
         aes_core_enc_block_n167, aes_core_enc_block_n166,
         aes_core_enc_block_n165, aes_core_enc_block_n164,
         aes_core_enc_block_n163, aes_core_enc_block_n162,
         aes_core_enc_block_n161, aes_core_enc_block_n160,
         aes_core_enc_block_n159, aes_core_enc_block_n158,
         aes_core_enc_block_n157, aes_core_enc_block_n156,
         aes_core_enc_block_n155, aes_core_enc_block_n154,
         aes_core_enc_block_n153, aes_core_enc_block_n152,
         aes_core_enc_block_n151, aes_core_enc_block_n150,
         aes_core_enc_block_n149, aes_core_enc_block_n148,
         aes_core_enc_block_n147, aes_core_enc_block_n146,
         aes_core_enc_block_n145, aes_core_enc_block_n144,
         aes_core_enc_block_n143, aes_core_enc_block_n142,
         aes_core_enc_block_n141, aes_core_enc_block_n140,
         aes_core_enc_block_n139, aes_core_enc_block_n138,
         aes_core_enc_block_n137, aes_core_enc_block_n136,
         aes_core_enc_block_n135, aes_core_enc_block_n134,
         aes_core_enc_block_n133, aes_core_enc_block_n132,
         aes_core_enc_block_n131, aes_core_enc_block_n130,
         aes_core_enc_block_n129, aes_core_enc_block_n128,
         aes_core_enc_block_n127, aes_core_enc_block_n126,
         aes_core_enc_block_n125, aes_core_enc_block_n124,
         aes_core_enc_block_n123, aes_core_enc_block_n122,
         aes_core_enc_block_n121, aes_core_enc_block_n120,
         aes_core_enc_block_n119, aes_core_enc_block_n118,
         aes_core_enc_block_n117, aes_core_enc_block_n116,
         aes_core_enc_block_n115, aes_core_enc_block_n114,
         aes_core_enc_block_n113, aes_core_enc_block_n112,
         aes_core_enc_block_n111, aes_core_enc_block_n110,
         aes_core_enc_block_n109, aes_core_enc_block_n108,
         aes_core_enc_block_n107, aes_core_enc_block_n106,
         aes_core_enc_block_n105, aes_core_enc_block_n104,
         aes_core_enc_block_n103, aes_core_enc_block_n102,
         aes_core_enc_block_n101, aes_core_enc_block_n100,
         aes_core_enc_block_n99, aes_core_enc_block_n98,
         aes_core_enc_block_n97, aes_core_enc_block_n96,
         aes_core_enc_block_n95, aes_core_enc_block_n94,
         aes_core_enc_block_n93, aes_core_enc_block_n92,
         aes_core_enc_block_n91, aes_core_enc_block_n90,
         aes_core_enc_block_n89, aes_core_enc_block_n88,
         aes_core_enc_block_n87, aes_core_enc_block_n86,
         aes_core_enc_block_n85, aes_core_enc_block_n84,
         aes_core_enc_block_n83, aes_core_enc_block_n82,
         aes_core_enc_block_n81, aes_core_enc_block_n80,
         aes_core_enc_block_n79, aes_core_enc_block_n78,
         aes_core_enc_block_n77, aes_core_enc_block_n76,
         aes_core_enc_block_n75, aes_core_enc_block_n74,
         aes_core_enc_block_n73, aes_core_enc_block_n72,
         aes_core_enc_block_n71, aes_core_enc_block_n70,
         aes_core_enc_block_n69, aes_core_enc_block_n68,
         aes_core_enc_block_n67, aes_core_enc_block_n66,
         aes_core_enc_block_n65, aes_core_enc_block_n64,
         aes_core_enc_block_n63, aes_core_enc_block_n62,
         aes_core_enc_block_n61, aes_core_enc_block_n60,
         aes_core_enc_block_n59, aes_core_enc_block_n58,
         aes_core_enc_block_n57, aes_core_enc_block_n56,
         aes_core_enc_block_n55, aes_core_enc_block_n54,
         aes_core_enc_block_n53, aes_core_enc_block_n52,
         aes_core_enc_block_n51, aes_core_enc_block_n50,
         aes_core_enc_block_n49, aes_core_enc_block_n48,
         aes_core_enc_block_n47, aes_core_enc_block_n46,
         aes_core_enc_block_n45, aes_core_enc_block_n44,
         aes_core_enc_block_n43, aes_core_enc_block_n42,
         aes_core_enc_block_n41, aes_core_enc_block_n40,
         aes_core_enc_block_n39, aes_core_enc_block_n38,
         aes_core_enc_block_n37, aes_core_enc_block_n36,
         aes_core_enc_block_n35, aes_core_enc_block_n34,
         aes_core_enc_block_n33, aes_core_enc_block_n32,
         aes_core_enc_block_n31, aes_core_enc_block_n30,
         aes_core_enc_block_n29, aes_core_enc_block_n28,
         aes_core_enc_block_n27, aes_core_enc_block_n26,
         aes_core_enc_block_n25, aes_core_enc_block_n24,
         aes_core_enc_block_n23, aes_core_enc_block_n22,
         aes_core_enc_block_n21, aes_core_enc_block_n20,
         aes_core_enc_block_n19, aes_core_enc_block_n18,
         aes_core_enc_block_n17, aes_core_enc_block_n16,
         aes_core_enc_block_n15, aes_core_enc_block_n14,
         aes_core_enc_block_n13, aes_core_enc_block_n12,
         aes_core_enc_block_n11, aes_core_enc_block_n10, aes_core_enc_block_n9,
         aes_core_enc_block_n8, aes_core_enc_block_n7, aes_core_enc_block_n6,
         aes_core_enc_block_n5, aes_core_enc_block_n4, aes_core_enc_block_n3,
         aes_core_enc_block_n2, aes_core_enc_block_n1,
         aes_core_enc_block_n1346, aes_core_enc_block_n1345,
         aes_core_enc_block_n1344, aes_core_enc_block_n1343,
         aes_core_enc_block_n1342, aes_core_enc_block_n1341,
         aes_core_enc_block_n1340, aes_core_enc_block_n1339,
         aes_core_enc_block_n1338, aes_core_enc_block_n1337,
         aes_core_enc_block_n1336, aes_core_enc_block_n1335,
         aes_core_enc_block_n1334, aes_core_enc_block_n1333,
         aes_core_enc_block_n1332, aes_core_enc_block_n1331,
         aes_core_enc_block_n1330, aes_core_enc_block_n1329,
         aes_core_enc_block_n1328, aes_core_enc_block_n1327,
         aes_core_enc_block_n1326, aes_core_enc_block_n1325,
         aes_core_enc_block_n1324, aes_core_enc_block_n1323,
         aes_core_enc_block_n1322, aes_core_enc_block_n1321,
         aes_core_enc_block_n1320, aes_core_enc_block_n1319,
         aes_core_enc_block_n1318, aes_core_enc_block_n1317,
         aes_core_enc_block_n1316, aes_core_enc_block_n1315,
         aes_core_enc_block_n1314, aes_core_enc_block_n1313,
         aes_core_enc_block_n1312, aes_core_enc_block_n1311,
         aes_core_enc_block_n1310, aes_core_enc_block_n1309,
         aes_core_enc_block_n1308, aes_core_enc_block_n1307,
         aes_core_enc_block_n1306, aes_core_enc_block_n1305,
         aes_core_enc_block_n1304, aes_core_enc_block_n1303,
         aes_core_enc_block_n1302, aes_core_enc_block_n1301,
         aes_core_enc_block_n1300, aes_core_enc_block_n1299,
         aes_core_enc_block_n1298, aes_core_enc_block_n1297,
         aes_core_enc_block_n1296, aes_core_enc_block_n1295,
         aes_core_enc_block_n1294, aes_core_enc_block_n1293,
         aes_core_enc_block_n1292, aes_core_enc_block_n1291,
         aes_core_enc_block_n1290, aes_core_enc_block_n1289,
         aes_core_enc_block_n1288, aes_core_enc_block_n1287,
         aes_core_enc_block_n1286, aes_core_enc_block_n1285,
         aes_core_enc_block_n1284, aes_core_enc_block_n1283,
         aes_core_enc_block_n1282, aes_core_enc_block_n1281,
         aes_core_enc_block_n1280, aes_core_enc_block_n1279,
         aes_core_enc_block_n1278, aes_core_enc_block_n1277,
         aes_core_enc_block_n1276, aes_core_enc_block_n1275,
         aes_core_enc_block_n1274, aes_core_enc_block_n1273,
         aes_core_enc_block_n1272, aes_core_enc_block_n1271,
         aes_core_enc_block_n1270, aes_core_enc_block_n1269,
         aes_core_enc_block_n1268, aes_core_enc_block_n1267,
         aes_core_enc_block_n1266, aes_core_enc_block_n1265,
         aes_core_enc_block_n1264, aes_core_enc_block_n1263,
         aes_core_enc_block_n1262, aes_core_enc_block_n1261,
         aes_core_enc_block_n1260, aes_core_enc_block_n1259,
         aes_core_enc_block_n1258, aes_core_enc_block_n1257,
         aes_core_enc_block_n1256, aes_core_enc_block_n1255,
         aes_core_enc_block_n1254, aes_core_enc_block_n1253,
         aes_core_enc_block_n1252, aes_core_enc_block_n1251,
         aes_core_enc_block_n1250, aes_core_enc_block_n1249,
         aes_core_enc_block_n1248, aes_core_enc_block_n1247,
         aes_core_enc_block_n1246, aes_core_enc_block_n1245,
         aes_core_enc_block_n1244, aes_core_enc_block_n1243,
         aes_core_enc_block_n1242, aes_core_enc_block_n1241,
         aes_core_enc_block_n1240, aes_core_enc_block_n1239,
         aes_core_enc_block_n1238, aes_core_enc_block_n1237,
         aes_core_enc_block_n1236, aes_core_enc_block_n1235,
         aes_core_enc_block_n1234, aes_core_enc_block_n1233,
         aes_core_enc_block_n1232, aes_core_enc_block_n1231,
         aes_core_enc_block_n1230, aes_core_enc_block_n1229,
         aes_core_enc_block_n1228, aes_core_enc_block_n1227,
         aes_core_enc_block_n1226, aes_core_enc_block_n1225,
         aes_core_enc_block_n1224, aes_core_enc_block_n1223,
         aes_core_enc_block_n1222, aes_core_enc_block_n1221,
         aes_core_enc_block_n1220, aes_core_enc_block_n1219,
         aes_core_enc_block_n1218, aes_core_enc_block_n1217,
         aes_core_enc_block_n1216, aes_core_enc_block_n1215,
         aes_core_enc_block_n1214, aes_core_enc_block_n1213,
         aes_core_enc_block_n1212, aes_core_enc_block_n1211,
         aes_core_enc_block_n1210, aes_core_enc_block_n1209,
         aes_core_enc_block_n1208, aes_core_enc_block_n1206,
         aes_core_enc_block_n1205, aes_core_enc_block_n1204,
         aes_core_enc_block_n1203, aes_core_enc_block_n1202,
         aes_core_enc_block_n1201, aes_core_enc_block_n1200,
         aes_core_enc_block_n1199, aes_core_enc_block_n1198,
         aes_core_enc_block_n1197, aes_core_enc_block_n1196,
         aes_core_enc_block_n1195, aes_core_enc_block_n1194,
         aes_core_enc_block_n1193, aes_core_enc_block_n1192,
         aes_core_enc_block_n1191, aes_core_enc_block_n1190,
         aes_core_enc_block_n1189, aes_core_enc_block_n1188,
         aes_core_enc_block_n1187, aes_core_enc_block_n1186,
         aes_core_enc_block_n1185, aes_core_enc_block_n1184,
         aes_core_enc_block_n1183, aes_core_enc_block_n1182,
         aes_core_enc_block_n1181, aes_core_enc_block_n1180,
         aes_core_enc_block_n1179, aes_core_enc_block_n1178,
         aes_core_enc_block_n1177, aes_core_enc_block_n1176,
         aes_core_enc_block_n1175, aes_core_enc_block_n1174,
         aes_core_enc_block_n1173, aes_core_enc_block_n1172,
         aes_core_enc_block_n1171, aes_core_enc_block_n1170,
         aes_core_enc_block_n1169, aes_core_enc_block_n1168,
         aes_core_enc_block_n1167, aes_core_enc_block_n1166,
         aes_core_enc_block_n1165, aes_core_enc_block_n1164,
         aes_core_enc_block_n1163, aes_core_enc_block_n1162,
         aes_core_enc_block_n1161, aes_core_enc_block_n1160,
         aes_core_enc_block_n1159, aes_core_enc_block_n1158,
         aes_core_enc_block_n1157, aes_core_enc_block_n1156,
         aes_core_enc_block_n1155, aes_core_enc_block_n1154,
         aes_core_enc_block_n1153, aes_core_enc_block_n1152,
         aes_core_enc_block_n1151, aes_core_enc_block_n1150,
         aes_core_enc_block_n1149, aes_core_enc_block_n1148,
         aes_core_enc_block_n1147, aes_core_enc_block_n1146,
         aes_core_enc_block_n1145, aes_core_enc_block_n1144,
         aes_core_enc_block_n1143, aes_core_enc_block_n1142,
         aes_core_enc_block_n1141, aes_core_enc_block_n1140,
         aes_core_enc_block_n1139, aes_core_enc_block_n1138,
         aes_core_enc_block_n1137, aes_core_enc_block_n1136,
         aes_core_enc_block_n1135, aes_core_enc_block_n1134,
         aes_core_enc_block_n1133, aes_core_enc_block_n1132,
         aes_core_enc_block_n1131, aes_core_enc_block_n1130,
         aes_core_enc_block_n1129, aes_core_enc_block_n1128,
         aes_core_enc_block_n1127, aes_core_enc_block_n1126,
         aes_core_enc_block_n1125, aes_core_enc_block_n1124,
         aes_core_enc_block_n1123, aes_core_enc_block_n1122,
         aes_core_enc_block_n1121, aes_core_enc_block_n1120,
         aes_core_enc_block_n1119, aes_core_enc_block_n1118,
         aes_core_enc_block_n1117, aes_core_enc_block_n1116,
         aes_core_enc_block_n1115, aes_core_enc_block_n1114,
         aes_core_enc_block_n1113, aes_core_enc_block_n1112,
         aes_core_enc_block_n1111, aes_core_enc_block_n1110,
         aes_core_enc_block_n1109, aes_core_enc_block_n1108,
         aes_core_enc_block_n1107, aes_core_enc_block_n1106,
         aes_core_enc_block_n1105, aes_core_enc_block_n1104,
         aes_core_enc_block_n1103, aes_core_enc_block_n1102,
         aes_core_enc_block_n1101, aes_core_enc_block_n1100,
         aes_core_enc_block_n1099, aes_core_enc_block_n1098,
         aes_core_enc_block_n1097, aes_core_enc_block_n1096,
         aes_core_enc_block_n1095, aes_core_enc_block_n1094,
         aes_core_enc_block_n1093, aes_core_enc_block_n1092,
         aes_core_enc_block_n1091, aes_core_enc_block_n1090,
         aes_core_enc_block_n1089, aes_core_enc_block_n1088,
         aes_core_enc_block_n1087, aes_core_enc_block_n1086,
         aes_core_enc_block_n1085, aes_core_enc_block_n1084,
         aes_core_enc_block_n1083, aes_core_enc_block_n1082,
         aes_core_enc_block_n1081, aes_core_enc_block_n1080,
         aes_core_enc_block_n1079, aes_core_enc_block_n1078,
         aes_core_enc_block_n1077, aes_core_enc_block_n1076,
         aes_core_enc_block_n1075, aes_core_enc_block_n1074,
         aes_core_enc_block_n1073, aes_core_enc_block_n1072,
         aes_core_enc_block_n1071, aes_core_enc_block_n1070,
         aes_core_enc_block_n1069, aes_core_enc_block_n1068,
         aes_core_enc_block_n1067, aes_core_enc_block_n1066,
         aes_core_enc_block_n1065, aes_core_enc_block_n1064,
         aes_core_enc_block_n1063, aes_core_enc_block_n1062,
         aes_core_enc_block_n1061, aes_core_enc_block_n1060,
         aes_core_enc_block_n1059, aes_core_enc_block_n1058,
         aes_core_enc_block_n1057, aes_core_enc_block_n1056,
         aes_core_enc_block_n1055, aes_core_enc_block_n1054,
         aes_core_enc_block_n1053, aes_core_enc_block_n1052,
         aes_core_enc_block_n1051, aes_core_enc_block_n1050,
         aes_core_enc_block_n1049, aes_core_enc_block_n1048,
         aes_core_enc_block_n1047, aes_core_enc_block_n1046,
         aes_core_enc_block_n1045, aes_core_enc_block_n1044,
         aes_core_enc_block_n1043, aes_core_enc_block_n1042,
         aes_core_enc_block_n1041, aes_core_enc_block_n1040,
         aes_core_enc_block_n1039, aes_core_enc_block_n1038,
         aes_core_enc_block_n1037, aes_core_enc_block_n1036,
         aes_core_enc_block_n1035, aes_core_enc_block_n1034,
         aes_core_enc_block_n1033, aes_core_enc_block_n1032,
         aes_core_enc_block_n1031, aes_core_enc_block_n1030,
         aes_core_enc_block_n1029, aes_core_enc_block_n1028,
         aes_core_enc_block_n1027, aes_core_enc_block_n1026,
         aes_core_enc_block_n1025, aes_core_enc_block_n1024,
         aes_core_enc_block_n1023, aes_core_enc_block_n1022,
         aes_core_enc_block_n1021, aes_core_enc_block_n1020,
         aes_core_enc_block_n1019, aes_core_enc_block_n1018,
         aes_core_enc_block_n1017, aes_core_enc_block_n1016,
         aes_core_enc_block_n1015, aes_core_enc_block_n1014,
         aes_core_enc_block_n1013, aes_core_enc_block_n1012,
         aes_core_enc_block_n1011, aes_core_enc_block_n1010,
         aes_core_enc_block_n1009, aes_core_enc_block_n1008,
         aes_core_enc_block_n1007, aes_core_enc_block_n1006,
         aes_core_enc_block_n1005, aes_core_enc_block_n1004,
         aes_core_enc_block_n1003, aes_core_enc_block_n1002,
         aes_core_enc_block_n1001, aes_core_enc_block_n1000,
         aes_core_enc_block_n999, aes_core_enc_block_n998,
         aes_core_enc_block_n997, aes_core_enc_block_n996,
         aes_core_enc_block_n995, aes_core_enc_block_n994,
         aes_core_enc_block_n993, aes_core_enc_block_n992,
         aes_core_enc_block_n991, aes_core_enc_block_n990,
         aes_core_enc_block_n989, aes_core_enc_block_n988,
         aes_core_enc_block_n987, aes_core_enc_block_n986,
         aes_core_enc_block_n985, aes_core_enc_block_n984,
         aes_core_enc_block_n983, aes_core_enc_block_n982,
         aes_core_enc_block_n981, aes_core_enc_block_n980,
         aes_core_enc_block_n979, aes_core_enc_block_n978,
         aes_core_enc_block_n977, aes_core_enc_block_n976,
         aes_core_enc_block_n975, aes_core_enc_block_n974,
         aes_core_enc_block_n973, aes_core_enc_block_n972,
         aes_core_enc_block_n971, aes_core_enc_block_n970,
         aes_core_enc_block_n969, aes_core_enc_block_n968,
         aes_core_enc_block_n967, aes_core_enc_block_n966,
         aes_core_enc_block_n965, aes_core_enc_block_n964,
         aes_core_enc_block_n963, aes_core_enc_block_n962,
         aes_core_enc_block_n961, aes_core_enc_block_n960,
         aes_core_enc_block_n959, aes_core_enc_block_n958,
         aes_core_enc_block_n957, aes_core_enc_block_n956,
         aes_core_enc_block_n955, aes_core_enc_block_n954,
         aes_core_enc_block_n953, aes_core_enc_block_n952,
         aes_core_enc_block_n951, aes_core_enc_block_n950,
         aes_core_enc_block_n949, aes_core_enc_block_n948,
         aes_core_enc_block_n946, aes_core_enc_block_n945,
         aes_core_enc_block_n944, aes_core_enc_block_n943,
         aes_core_enc_block_n942, aes_core_enc_block_n941,
         aes_core_enc_block_n940, aes_core_enc_block_n939,
         aes_core_enc_block_n938, aes_core_enc_block_n937,
         aes_core_enc_block_n936, aes_core_enc_block_n935,
         aes_core_enc_block_n934, aes_core_enc_block_n933,
         aes_core_enc_block_n932, aes_core_enc_block_n931,
         aes_core_enc_block_n930, aes_core_enc_block_n929,
         aes_core_enc_block_n928, aes_core_enc_block_n927,
         aes_core_enc_block_n926, aes_core_enc_block_n925,
         aes_core_enc_block_n924, aes_core_enc_block_n923,
         aes_core_enc_block_n922, aes_core_enc_block_n921,
         aes_core_enc_block_n920, aes_core_enc_block_n919,
         aes_core_enc_block_n918, aes_core_enc_block_n917,
         aes_core_enc_block_n916, aes_core_enc_block_n915,
         aes_core_enc_block_n914, aes_core_enc_block_n913,
         aes_core_enc_block_n912, aes_core_enc_block_n911,
         aes_core_enc_block_n910, aes_core_enc_block_n909,
         aes_core_enc_block_n908, aes_core_enc_block_n907,
         aes_core_enc_block_n906, aes_core_enc_block_n905,
         aes_core_enc_block_n904, aes_core_enc_block_n903,
         aes_core_enc_block_n902, aes_core_enc_block_n901,
         aes_core_enc_block_n900, aes_core_enc_block_n899,
         aes_core_enc_block_n898, aes_core_enc_block_n897,
         aes_core_enc_block_n896, aes_core_enc_block_n895,
         aes_core_enc_block_n894, aes_core_enc_block_n893,
         aes_core_enc_block_n892, aes_core_enc_block_n891,
         aes_core_enc_block_n890, aes_core_enc_block_n889,
         aes_core_enc_block_n888, aes_core_enc_block_n887,
         aes_core_enc_block_n886, aes_core_enc_block_n885,
         aes_core_enc_block_n884, aes_core_enc_block_n883,
         aes_core_enc_block_n882, aes_core_enc_block_n881,
         aes_core_enc_block_n880, aes_core_enc_block_n879,
         aes_core_enc_block_n878, aes_core_enc_block_n877,
         aes_core_enc_block_n876, aes_core_enc_block_n875,
         aes_core_enc_block_n874, aes_core_enc_block_n873,
         aes_core_enc_block_n872, aes_core_enc_block_n871,
         aes_core_enc_block_n870, aes_core_enc_block_n869,
         aes_core_enc_block_n868, aes_core_enc_block_n867,
         aes_core_enc_block_n866, aes_core_enc_block_n865,
         aes_core_enc_block_n864, aes_core_enc_block_n863,
         aes_core_enc_block_n862, aes_core_enc_block_n861,
         aes_core_enc_block_n860, aes_core_enc_block_n859,
         aes_core_enc_block_n858, aes_core_enc_block_n857,
         aes_core_enc_block_n856, aes_core_enc_block_n855,
         aes_core_enc_block_n854, aes_core_enc_block_n853,
         aes_core_enc_block_n852, aes_core_enc_block_n851,
         aes_core_enc_block_n850, aes_core_enc_block_n849,
         aes_core_enc_block_n848, aes_core_enc_block_n847,
         aes_core_enc_block_n846, aes_core_enc_block_n845,
         aes_core_enc_block_n844, aes_core_enc_block_n843,
         aes_core_enc_block_n842, aes_core_enc_block_n841,
         aes_core_enc_block_n840, aes_core_enc_block_n839,
         aes_core_enc_block_n838, aes_core_enc_block_n837,
         aes_core_enc_block_n836, aes_core_enc_block_n835,
         aes_core_enc_block_n834, aes_core_enc_block_n833,
         aes_core_enc_block_n832, aes_core_enc_block_n831,
         aes_core_enc_block_n830, aes_core_enc_block_n829,
         aes_core_enc_block_n828, aes_core_enc_block_n827,
         aes_core_enc_block_n826, aes_core_enc_block_n825,
         aes_core_enc_block_n824, aes_core_enc_block_n823,
         aes_core_enc_block_n822, aes_core_enc_block_n821,
         aes_core_enc_block_n820, aes_core_enc_block_n819,
         aes_core_enc_block_n818, aes_core_enc_block_n817,
         aes_core_enc_block_n816, aes_core_enc_block_n815,
         aes_core_enc_block_n814, aes_core_enc_block_n813,
         aes_core_enc_block_n812, aes_core_enc_block_n811,
         aes_core_enc_block_n810, aes_core_enc_block_n809,
         aes_core_enc_block_n808, aes_core_enc_block_n807,
         aes_core_enc_block_n806, aes_core_enc_block_n805,
         aes_core_enc_block_n804, aes_core_enc_block_n803,
         aes_core_enc_block_n802, aes_core_enc_block_n801,
         aes_core_enc_block_n800, aes_core_enc_block_n799,
         aes_core_enc_block_n798, aes_core_enc_block_n797,
         aes_core_enc_block_n796, aes_core_enc_block_n795,
         aes_core_enc_block_n794, aes_core_enc_block_n793,
         aes_core_enc_block_n792, aes_core_enc_block_n791,
         aes_core_enc_block_n790, aes_core_enc_block_n789,
         aes_core_enc_block_n788, aes_core_enc_block_n787,
         aes_core_enc_block_n786, aes_core_enc_block_n785,
         aes_core_enc_block_n784, aes_core_enc_block_n783,
         aes_core_enc_block_n782, aes_core_enc_block_n781,
         aes_core_enc_block_n780, aes_core_enc_block_n779,
         aes_core_enc_block_n778, aes_core_enc_block_n777,
         aes_core_enc_block_n776, aes_core_enc_block_n775,
         aes_core_enc_block_n774, aes_core_enc_block_n773,
         aes_core_enc_block_n772, aes_core_enc_block_n771,
         aes_core_enc_block_n770, aes_core_enc_block_n769,
         aes_core_enc_block_n768, aes_core_enc_block_n767,
         aes_core_enc_block_n766, aes_core_enc_block_n765,
         aes_core_enc_block_n764, aes_core_enc_block_n763,
         aes_core_enc_block_n762, aes_core_enc_block_n761,
         aes_core_enc_block_n760, aes_core_enc_block_n759,
         aes_core_enc_block_n758, aes_core_enc_block_n757,
         aes_core_enc_block_n756, aes_core_enc_block_n755,
         aes_core_enc_block_n754, aes_core_enc_block_n753,
         aes_core_enc_block_n752, aes_core_enc_block_n751,
         aes_core_enc_block_n750, aes_core_enc_block_n749,
         aes_core_enc_block_n748, aes_core_enc_block_n747,
         aes_core_enc_block_n746, aes_core_enc_block_n745,
         aes_core_enc_block_n744, aes_core_enc_block_n743,
         aes_core_enc_block_n742, aes_core_enc_block_n741,
         aes_core_enc_block_n740, aes_core_enc_block_n739,
         aes_core_enc_block_n738, aes_core_enc_block_n737,
         aes_core_enc_block_n736, aes_core_enc_block_n735,
         aes_core_enc_block_n734, aes_core_enc_block_n733,
         aes_core_enc_block_n732, aes_core_enc_block_n731,
         aes_core_enc_block_n730, aes_core_enc_block_n729,
         aes_core_enc_block_n728, aes_core_enc_block_n727,
         aes_core_enc_block_n726, aes_core_enc_block_n725,
         aes_core_enc_block_n724, aes_core_enc_block_n723,
         aes_core_enc_block_n722, aes_core_enc_block_n721,
         aes_core_enc_block_n720, aes_core_enc_block_n719,
         aes_core_enc_block_n718, aes_core_enc_block_n717,
         aes_core_enc_block_n716, aes_core_enc_block_n715,
         aes_core_enc_block_n714, aes_core_enc_block_n713,
         aes_core_enc_block_n712, aes_core_enc_block_n711,
         aes_core_enc_block_n710, aes_core_enc_block_n709,
         aes_core_enc_block_n707, aes_core_enc_block_n706,
         aes_core_enc_block_n705, aes_core_enc_block_n704,
         aes_core_enc_block_n703, aes_core_enc_block_n702,
         aes_core_enc_block_n701, aes_core_enc_block_n700,
         aes_core_enc_block_n699, aes_core_enc_block_n698,
         aes_core_enc_block_n697, aes_core_enc_block_n696,
         aes_core_enc_block_n695, aes_core_enc_block_n694,
         aes_core_enc_block_n693, aes_core_enc_block_n692,
         aes_core_enc_block_n691, aes_core_enc_block_n690,
         aes_core_enc_block_n689, aes_core_enc_block_n688,
         aes_core_enc_block_n687, aes_core_enc_block_n686,
         aes_core_enc_block_n685, aes_core_enc_block_n684,
         aes_core_enc_block_n683, aes_core_enc_block_n682,
         aes_core_enc_block_n681, aes_core_enc_block_n680,
         aes_core_enc_block_n679, aes_core_enc_block_n678,
         aes_core_enc_block_n677, aes_core_enc_block_n676,
         aes_core_enc_block_n675, aes_core_enc_block_n674,
         aes_core_enc_block_n673, aes_core_enc_block_n672,
         aes_core_enc_block_n671, aes_core_enc_block_n670,
         aes_core_enc_block_n669, aes_core_enc_block_n668,
         aes_core_enc_block_n667, aes_core_enc_block_n666,
         aes_core_enc_block_n665, aes_core_enc_block_n664,
         aes_core_enc_block_n663, aes_core_enc_block_n662,
         aes_core_enc_block_n661, aes_core_enc_block_n660,
         aes_core_enc_block_n659, aes_core_enc_block_n658,
         aes_core_enc_block_n657, aes_core_enc_block_n656,
         aes_core_enc_block_n655, aes_core_enc_block_n654,
         aes_core_enc_block_n653, aes_core_enc_block_n652,
         aes_core_enc_block_n651, aes_core_enc_block_n650,
         aes_core_enc_block_n649, aes_core_enc_block_n648,
         aes_core_enc_block_n647, aes_core_enc_block_n646,
         aes_core_enc_block_n645, aes_core_enc_block_n644,
         aes_core_enc_block_n643, aes_core_enc_block_n642,
         aes_core_enc_block_n641, aes_core_enc_block_n640,
         aes_core_enc_block_n639, aes_core_enc_block_n638,
         aes_core_enc_block_n637, aes_core_enc_block_n636,
         aes_core_enc_block_n635, aes_core_enc_block_n634,
         aes_core_enc_block_n633, aes_core_enc_block_n632,
         aes_core_enc_block_n631, aes_core_enc_block_n630,
         aes_core_enc_block_n629, aes_core_enc_block_n628,
         aes_core_enc_block_n627, aes_core_enc_block_n626,
         aes_core_enc_block_n625, aes_core_enc_block_n624,
         aes_core_enc_block_n623, aes_core_enc_block_n622,
         aes_core_enc_block_n621, aes_core_enc_block_n620,
         aes_core_enc_block_n619, aes_core_enc_block_n618,
         aes_core_enc_block_n617, aes_core_enc_block_n616,
         aes_core_enc_block_n615, aes_core_enc_block_n614,
         aes_core_enc_block_n613, aes_core_enc_block_n612,
         aes_core_enc_block_n611, aes_core_enc_block_n610,
         aes_core_enc_block_n609, aes_core_enc_block_n608,
         aes_core_enc_block_n607, aes_core_enc_block_n606,
         aes_core_enc_block_n605, aes_core_enc_block_n604,
         aes_core_enc_block_n603, aes_core_enc_block_n602,
         aes_core_enc_block_n601, aes_core_enc_block_n600,
         aes_core_enc_block_n599, aes_core_enc_block_n598,
         aes_core_enc_block_n597, aes_core_enc_block_n596,
         aes_core_enc_block_n595, aes_core_enc_block_n594,
         aes_core_enc_block_n593, aes_core_enc_block_n592,
         aes_core_enc_block_n591, aes_core_enc_block_n590,
         aes_core_enc_block_n589, aes_core_enc_block_n588,
         aes_core_enc_block_n587, aes_core_enc_block_n586,
         aes_core_enc_block_n585, aes_core_enc_block_n584,
         aes_core_enc_block_n583, aes_core_enc_block_n582,
         aes_core_enc_block_n581, aes_core_enc_block_n580,
         aes_core_enc_block_n579, aes_core_enc_block_n578,
         aes_core_enc_block_n577, aes_core_enc_block_n576,
         aes_core_enc_block_n575, aes_core_enc_block_n574,
         aes_core_enc_block_n573, aes_core_enc_block_n572,
         aes_core_enc_block_n571, aes_core_enc_block_n570,
         aes_core_enc_block_n569, aes_core_enc_block_n568,
         aes_core_enc_block_n567, aes_core_enc_block_n566,
         aes_core_enc_block_n565, aes_core_enc_block_n564,
         aes_core_enc_block_n563, aes_core_enc_block_n562,
         aes_core_enc_block_n561, aes_core_enc_block_n560,
         aes_core_enc_block_n559, aes_core_enc_block_n558,
         aes_core_enc_block_n557, aes_core_enc_block_n556,
         aes_core_enc_block_n555, aes_core_enc_block_n554,
         aes_core_enc_block_n553, aes_core_enc_block_n552,
         aes_core_enc_block_n551, aes_core_enc_block_n550,
         aes_core_enc_block_n549, aes_core_enc_block_n548,
         aes_core_enc_block_n547, aes_core_enc_block_n546,
         aes_core_enc_block_n545, aes_core_enc_block_n544,
         aes_core_enc_block_n543, aes_core_enc_block_n542,
         aes_core_enc_block_n541, aes_core_enc_block_n540,
         aes_core_enc_block_n539, aes_core_enc_block_n538,
         aes_core_enc_block_n537, aes_core_enc_block_n536,
         aes_core_enc_block_n535, aes_core_enc_block_n534,
         aes_core_enc_block_n533, aes_core_enc_block_n532,
         aes_core_enc_block_n531, aes_core_enc_block_n530,
         aes_core_enc_block_n529, aes_core_enc_block_n528,
         aes_core_enc_block_n527, aes_core_enc_block_n526,
         aes_core_enc_block_n525, aes_core_enc_block_n524,
         aes_core_enc_block_n523, aes_core_enc_block_n522,
         aes_core_enc_block_n521, aes_core_enc_block_n520,
         aes_core_enc_block_n519, aes_core_enc_block_n518,
         aes_core_enc_block_n517, aes_core_enc_block_n516,
         aes_core_enc_block_n515, aes_core_enc_block_n514,
         aes_core_enc_block_n513, aes_core_enc_block_n512,
         aes_core_enc_block_n511, aes_core_enc_block_n510,
         aes_core_enc_block_n509, aes_core_enc_block_n508,
         aes_core_enc_block_n507, aes_core_enc_block_n506,
         aes_core_enc_block_n505, aes_core_enc_block_n504,
         aes_core_enc_block_n503, aes_core_enc_block_n502,
         aes_core_enc_block_n501, aes_core_enc_block_n500,
         aes_core_enc_block_n499, aes_core_enc_block_n498,
         aes_core_enc_block_n497, aes_core_enc_block_n496,
         aes_core_enc_block_n495, aes_core_enc_block_n494,
         aes_core_enc_block_n493, aes_core_enc_block_n492,
         aes_core_enc_block_n491, aes_core_enc_block_n490,
         aes_core_enc_block_n489, aes_core_enc_block_n488,
         aes_core_enc_block_n487, aes_core_enc_block_n486,
         aes_core_enc_block_n485, aes_core_enc_block_n484,
         aes_core_enc_block_n483, aes_core_enc_block_n482,
         aes_core_enc_block_n481, aes_core_enc_block_n480,
         aes_core_enc_block_n479, aes_core_enc_block_n478,
         aes_core_enc_block_n477, aes_core_enc_block_n476,
         aes_core_enc_block_n475, aes_core_enc_block_n474,
         aes_core_enc_block_n473, aes_core_enc_block_n472,
         aes_core_enc_block_n471, aes_core_enc_block_n470,
         aes_core_enc_block_n469, aes_core_enc_block_n468,
         aes_core_enc_block_n466, aes_core_enc_block_n465,
         aes_core_enc_block_n464, aes_core_enc_block_n463,
         aes_core_enc_block_n462, aes_core_enc_block_n461,
         aes_core_enc_block_n460, aes_core_enc_block_n459,
         aes_core_enc_block_n458, aes_core_enc_block_n457,
         aes_core_enc_block_n456, aes_core_enc_block_n455,
         aes_core_enc_block_n454, aes_core_enc_block_n453,
         aes_core_enc_block_n452, aes_core_enc_block_n451,
         aes_core_enc_block_n450, aes_core_enc_block_n449,
         aes_core_enc_block_n448, aes_core_enc_block_n447,
         aes_core_enc_block_n446, aes_core_enc_block_n445,
         aes_core_enc_block_n444, aes_core_enc_block_n443,
         aes_core_enc_block_n442, aes_core_enc_block_n441,
         aes_core_enc_block_n440, aes_core_enc_block_n439,
         aes_core_enc_block_n438, aes_core_enc_block_n437,
         aes_core_enc_block_n436, aes_core_enc_block_n435,
         aes_core_enc_block_n434, aes_core_enc_block_n433,
         aes_core_enc_block_n432, aes_core_enc_block_n431,
         aes_core_enc_block_n430, aes_core_enc_block_n429,
         aes_core_enc_block_n428, aes_core_enc_block_n427,
         aes_core_enc_block_n426, aes_core_enc_block_n425,
         aes_core_enc_block_n424, aes_core_enc_block_n423,
         aes_core_enc_block_n422, aes_core_enc_block_n421,
         aes_core_enc_block_n420, aes_core_enc_block_n419,
         aes_core_enc_block_n418, aes_core_enc_block_n417,
         aes_core_enc_block_n416, aes_core_enc_block_n415,
         aes_core_enc_block_n414, aes_core_enc_block_n413,
         aes_core_enc_block_n412, aes_core_enc_block_n411,
         aes_core_enc_block_n410, aes_core_enc_block_n409,
         aes_core_enc_block_n408, aes_core_enc_block_n407,
         aes_core_enc_block_n406, aes_core_enc_block_n405,
         aes_core_enc_block_n404, aes_core_enc_block_n403,
         aes_core_enc_block_n402, aes_core_enc_block_n401,
         aes_core_enc_block_n400, aes_core_enc_block_n399,
         aes_core_enc_block_n398, aes_core_enc_block_n397,
         aes_core_enc_block_n396, aes_core_enc_block_n395,
         aes_core_enc_block_n394, aes_core_enc_block_n393,
         aes_core_enc_block_n392, aes_core_enc_block_n391,
         aes_core_enc_block_n390, aes_core_enc_block_n389,
         aes_core_enc_block_n388, aes_core_enc_block_n387,
         aes_core_enc_block_n386, aes_core_enc_block_n385,
         aes_core_enc_block_n384, aes_core_enc_block_n383,
         aes_core_enc_block_n382, aes_core_enc_block_n381,
         aes_core_enc_block_n380, aes_core_enc_block_n379,
         aes_core_enc_block_n378, aes_core_enc_block_n377,
         aes_core_enc_block_n376, aes_core_enc_block_n375,
         aes_core_enc_block_n374, aes_core_enc_block_n373,
         aes_core_enc_block_n372, aes_core_enc_block_n371,
         aes_core_enc_block_n370, aes_core_enc_block_n369,
         aes_core_enc_block_n368, aes_core_enc_block_n367,
         aes_core_enc_block_n366, aes_core_enc_block_n365,
         aes_core_enc_block_n364, aes_core_enc_block_n363,
         aes_core_enc_block_n362, aes_core_enc_block_n361,
         aes_core_enc_block_n360, aes_core_enc_block_n359,
         aes_core_enc_block_n358, aes_core_enc_block_n357,
         aes_core_enc_block_n356, aes_core_enc_block_n355,
         aes_core_enc_block_n354, aes_core_enc_block_n353,
         aes_core_enc_block_n352, aes_core_enc_block_n351,
         aes_core_enc_block_n350, aes_core_enc_block_n349,
         aes_core_enc_block_n348, aes_core_enc_block_n347,
         aes_core_enc_block_n346, aes_core_enc_block_n345,
         aes_core_enc_block_n344, aes_core_enc_block_n343,
         aes_core_enc_block_n342, aes_core_enc_block_n341,
         aes_core_enc_block_n340, aes_core_enc_block_n339,
         aes_core_enc_block_n338, aes_core_enc_block_n337,
         aes_core_enc_block_n336, aes_core_enc_block_n335,
         aes_core_enc_block_n334, aes_core_enc_block_n333,
         aes_core_enc_block_n332, aes_core_enc_block_n331,
         aes_core_enc_block_n330, aes_core_enc_block_n329,
         aes_core_enc_block_n328, aes_core_enc_block_n327,
         aes_core_enc_block_n326, aes_core_enc_block_n325,
         aes_core_enc_block_n324, aes_core_enc_block_n323,
         aes_core_enc_block_n322, aes_core_enc_block_n321,
         aes_core_enc_block_n320, aes_core_enc_block_n319,
         aes_core_enc_block_n318, aes_core_enc_block_n317,
         aes_core_enc_block_n316, aes_core_enc_block_n315,
         aes_core_enc_block_n314, aes_core_enc_block_n313,
         aes_core_enc_block_n312, aes_core_enc_block_n311,
         aes_core_enc_block_n310, aes_core_enc_block_n309,
         aes_core_enc_block_n308, aes_core_enc_block_n307,
         aes_core_enc_block_n306, aes_core_enc_block_n305,
         aes_core_enc_block_n304, aes_core_enc_block_n303,
         aes_core_enc_block_n302, aes_core_enc_block_n301,
         aes_core_enc_block_n300, aes_core_enc_block_n299,
         aes_core_enc_block_n298, aes_core_enc_block_n297,
         aes_core_enc_block_n296, aes_core_enc_block_n295,
         aes_core_enc_block_n294, aes_core_enc_block_n293,
         aes_core_enc_block_n292, aes_core_enc_block_n291,
         aes_core_enc_block_n290, aes_core_enc_block_n289,
         aes_core_enc_block_n288, aes_core_enc_block_n287,
         aes_core_enc_block_n286, aes_core_enc_block_n285,
         aes_core_enc_block_n284, aes_core_enc_block_n283,
         aes_core_enc_block_n282, aes_core_enc_block_n281,
         aes_core_enc_block_n280, aes_core_enc_block_n279,
         aes_core_enc_block_n278, aes_core_enc_block_n277,
         aes_core_enc_block_n276, aes_core_enc_block_n275,
         aes_core_enc_block_n274, aes_core_enc_block_n273,
         aes_core_enc_block_n272, aes_core_enc_block_n271,
         aes_core_enc_block_n270, aes_core_enc_block_n269,
         aes_core_enc_block_n268, aes_core_enc_block_n267,
         aes_core_enc_block_n266, aes_core_enc_block_n265,
         aes_core_enc_block_n264, aes_core_enc_block_n263,
         aes_core_enc_block_n262, aes_core_enc_block_n261,
         aes_core_enc_block_n260, aes_core_enc_block_n259,
         aes_core_enc_block_n258, aes_core_enc_block_n257,
         aes_core_enc_block_n256, aes_core_enc_block_n255,
         aes_core_enc_block_n254, aes_core_enc_block_n253,
         aes_core_enc_block_n252, aes_core_enc_block_n251,
         aes_core_enc_block_n250, aes_core_enc_block_n249,
         aes_core_enc_block_n248, aes_core_enc_block_n247,
         aes_core_enc_block_n246, aes_core_enc_block_n245,
         aes_core_enc_block_n244, aes_core_enc_block_n243,
         aes_core_enc_block_n242, aes_core_enc_block_n241,
         aes_core_enc_block_n239, aes_core_enc_block_n238,
         aes_core_enc_block_n237, aes_core_enc_block_n236,
         aes_core_enc_block_n235, aes_core_enc_block_n234,
         aes_core_enc_block_n233, aes_core_enc_block_n231,
         aes_core_enc_block_n230, aes_core_enc_block_n229,
         aes_core_enc_block_n228, aes_core_enc_block_n227,
         aes_core_enc_block_n226, aes_core_enc_block_n225,
         aes_core_enc_block_n224, aes_core_enc_block_n223,
         aes_core_enc_block_n222, aes_core_enc_block_n221,
         aes_core_enc_block_n220, aes_core_enc_block_n219,
         aes_core_enc_block_n218, aes_core_enc_block_n217,
         aes_core_enc_block_n216, aes_core_enc_block_n215,
         aes_core_enc_block_n214, aes_core_enc_block_n213,
         aes_core_enc_block_n212, aes_core_enc_block_n211,
         aes_core_enc_block_n210, aes_core_enc_block_n209,
         aes_core_enc_block_n208, aes_core_enc_block_n207,
         aes_core_enc_block_n206, aes_core_enc_block_n205,
         aes_core_enc_block_n204, aes_core_enc_block_n203,
         aes_core_enc_block_n202, aes_core_enc_block_n201,
         aes_core_enc_block_n200, aes_core_enc_block_n199,
         aes_core_enc_block_n198, aes_core_enc_block_n197,
         aes_core_keymem_n2773, aes_core_keymem_n2772, aes_core_keymem_n2771,
         aes_core_keymem_n2770, aes_core_keymem_n2769, aes_core_keymem_n2768,
         aes_core_keymem_n2767, aes_core_keymem_n2766, aes_core_keymem_n2765,
         aes_core_keymem_n2764, aes_core_keymem_n2763, aes_core_keymem_n2762,
         aes_core_keymem_n2761, aes_core_keymem_n2760, aes_core_keymem_n2759,
         aes_core_keymem_n2758, aes_core_keymem_n2757, aes_core_keymem_n2756,
         aes_core_keymem_n2755, aes_core_keymem_n2754, aes_core_keymem_n2753,
         aes_core_keymem_n2752, aes_core_keymem_n2751, aes_core_keymem_n2750,
         aes_core_keymem_n2749, aes_core_keymem_n2748, aes_core_keymem_n2747,
         aes_core_keymem_n2746, aes_core_keymem_n2745, aes_core_keymem_n2744,
         aes_core_keymem_n2743, aes_core_keymem_n2742, aes_core_keymem_n2741,
         aes_core_keymem_n2740, aes_core_keymem_n2739, aes_core_keymem_n2738,
         aes_core_keymem_n2737, aes_core_keymem_n2736, aes_core_keymem_n2735,
         aes_core_keymem_n2734, aes_core_keymem_n2733, aes_core_keymem_n2732,
         aes_core_keymem_n2731, aes_core_keymem_n2730, aes_core_keymem_n2729,
         aes_core_keymem_n2728, aes_core_keymem_n2727, aes_core_keymem_n2726,
         aes_core_keymem_n2725, aes_core_keymem_n2724, aes_core_keymem_n2723,
         aes_core_keymem_n2722, aes_core_keymem_n2721, aes_core_keymem_n2720,
         aes_core_keymem_n2719, aes_core_keymem_n2718, aes_core_keymem_n2717,
         aes_core_keymem_n2716, aes_core_keymem_n2715, aes_core_keymem_n2714,
         aes_core_keymem_n2713, aes_core_keymem_n2712, aes_core_keymem_n2711,
         aes_core_keymem_n2710, aes_core_keymem_n2709, aes_core_keymem_n2708,
         aes_core_keymem_n2707, aes_core_keymem_n2706, aes_core_keymem_n2705,
         aes_core_keymem_n2704, aes_core_keymem_n2703, aes_core_keymem_n2702,
         aes_core_keymem_n2701, aes_core_keymem_n2700, aes_core_keymem_n2699,
         aes_core_keymem_n2698, aes_core_keymem_n2697, aes_core_keymem_n2696,
         aes_core_keymem_n2695, aes_core_keymem_n2694, aes_core_keymem_n2693,
         aes_core_keymem_n2692, aes_core_keymem_n2691, aes_core_keymem_n2690,
         aes_core_keymem_n2689, aes_core_keymem_n2688, aes_core_keymem_n2687,
         aes_core_keymem_n2686, aes_core_keymem_n2685, aes_core_keymem_n2684,
         aes_core_keymem_n2683, aes_core_keymem_n2682, aes_core_keymem_n2681,
         aes_core_keymem_n2680, aes_core_keymem_n2679, aes_core_keymem_n2678,
         aes_core_keymem_n2677, aes_core_keymem_n2676, aes_core_keymem_n2675,
         aes_core_keymem_n2674, aes_core_keymem_n2673, aes_core_keymem_n2672,
         aes_core_keymem_n2671, aes_core_keymem_n2670, aes_core_keymem_n2669,
         aes_core_keymem_n2668, aes_core_keymem_n2667, aes_core_keymem_n2666,
         aes_core_keymem_n2665, aes_core_keymem_n2664, aes_core_keymem_n2663,
         aes_core_keymem_n2662, aes_core_keymem_n2661, aes_core_keymem_n2660,
         aes_core_keymem_n2659, aes_core_keymem_n2658, aes_core_keymem_n2657,
         aes_core_keymem_n2656, aes_core_keymem_n2655, aes_core_keymem_n2654,
         aes_core_keymem_n2653, aes_core_keymem_n2652, aes_core_keymem_n2651,
         aes_core_keymem_n2650, aes_core_keymem_n2649, aes_core_keymem_n2648,
         aes_core_keymem_n2647, aes_core_keymem_n2646, aes_core_keymem_n2645,
         aes_core_keymem_n2644, aes_core_keymem_n2643, aes_core_keymem_n2642,
         aes_core_keymem_n2641, aes_core_keymem_n2640, aes_core_keymem_n2639,
         aes_core_keymem_n2638, aes_core_keymem_n2637, aes_core_keymem_n2636,
         aes_core_keymem_n2635, aes_core_keymem_n2634, aes_core_keymem_n2633,
         aes_core_keymem_n2632, aes_core_keymem_n2631, aes_core_keymem_n2630,
         aes_core_keymem_n2629, aes_core_keymem_n2628, aes_core_keymem_n2627,
         aes_core_keymem_n2626, aes_core_keymem_n2625, aes_core_keymem_n2624,
         aes_core_keymem_n2623, aes_core_keymem_n2622, aes_core_keymem_n2621,
         aes_core_keymem_n2620, aes_core_keymem_n2619, aes_core_keymem_n2618,
         aes_core_keymem_n2617, aes_core_keymem_n2616, aes_core_keymem_n2615,
         aes_core_keymem_n2614, aes_core_keymem_n2613, aes_core_keymem_n2612,
         aes_core_keymem_n2611, aes_core_keymem_n2610, aes_core_keymem_n2609,
         aes_core_keymem_n2608, aes_core_keymem_n2607, aes_core_keymem_n2606,
         aes_core_keymem_n2605, aes_core_keymem_n2604, aes_core_keymem_n2603,
         aes_core_keymem_n2602, aes_core_keymem_n2601, aes_core_keymem_n2600,
         aes_core_keymem_n2599, aes_core_keymem_n2598, aes_core_keymem_n2597,
         aes_core_keymem_n2596, aes_core_keymem_n2595, aes_core_keymem_n2594,
         aes_core_keymem_n2593, aes_core_keymem_n2592, aes_core_keymem_n2591,
         aes_core_keymem_n2590, aes_core_keymem_n2589, aes_core_keymem_n2588,
         aes_core_keymem_n2587, aes_core_keymem_n2586, aes_core_keymem_n2585,
         aes_core_keymem_n2584, aes_core_keymem_n2583, aes_core_keymem_n2582,
         aes_core_keymem_n2581, aes_core_keymem_n2580, aes_core_keymem_n2579,
         aes_core_keymem_n2578, aes_core_keymem_n2577, aes_core_keymem_n2576,
         aes_core_keymem_n2575, aes_core_keymem_n2574, aes_core_keymem_n2573,
         aes_core_keymem_n2572, aes_core_keymem_n2571, aes_core_keymem_n2570,
         aes_core_keymem_n2569, aes_core_keymem_n2568, aes_core_keymem_n2567,
         aes_core_keymem_n2566, aes_core_keymem_n2565, aes_core_keymem_n2564,
         aes_core_keymem_n2563, aes_core_keymem_n2562, aes_core_keymem_n2561,
         aes_core_keymem_n2560, aes_core_keymem_n2559, aes_core_keymem_n2558,
         aes_core_keymem_n2557, aes_core_keymem_n2556, aes_core_keymem_n2555,
         aes_core_keymem_n2554, aes_core_keymem_n2553, aes_core_keymem_n2552,
         aes_core_keymem_n2551, aes_core_keymem_n2550, aes_core_keymem_n2549,
         aes_core_keymem_n2548, aes_core_keymem_n2547, aes_core_keymem_n2546,
         aes_core_keymem_n2545, aes_core_keymem_n2544, aes_core_keymem_n2543,
         aes_core_keymem_n2542, aes_core_keymem_n2541, aes_core_keymem_n2540,
         aes_core_keymem_n2539, aes_core_keymem_n2538, aes_core_keymem_n2537,
         aes_core_keymem_n2536, aes_core_keymem_n2535, aes_core_keymem_n2534,
         aes_core_keymem_n2533, aes_core_keymem_n2532, aes_core_keymem_n2531,
         aes_core_keymem_n2530, aes_core_keymem_n2529, aes_core_keymem_n2528,
         aes_core_keymem_n2527, aes_core_keymem_n2526, aes_core_keymem_n2525,
         aes_core_keymem_n2524, aes_core_keymem_n2523, aes_core_keymem_n2522,
         aes_core_keymem_n2521, aes_core_keymem_n2520, aes_core_keymem_n2519,
         aes_core_keymem_n2518, aes_core_keymem_n2517, aes_core_keymem_n2516,
         aes_core_keymem_n2515, aes_core_keymem_n2514, aes_core_keymem_n2513,
         aes_core_keymem_n2512, aes_core_keymem_n2511, aes_core_keymem_n2510,
         aes_core_keymem_n2509, aes_core_keymem_n2508, aes_core_keymem_n2507,
         aes_core_keymem_n2506, aes_core_keymem_n2505, aes_core_keymem_n2504,
         aes_core_keymem_n2503, aes_core_keymem_n2502, aes_core_keymem_n2501,
         aes_core_keymem_n2500, aes_core_keymem_n2499, aes_core_keymem_n2498,
         aes_core_keymem_n2497, aes_core_keymem_n2496, aes_core_keymem_n2495,
         aes_core_keymem_n2494, aes_core_keymem_n2493, aes_core_keymem_n2492,
         aes_core_keymem_n2491, aes_core_keymem_n2490, aes_core_keymem_n2489,
         aes_core_keymem_n2488, aes_core_keymem_n2487, aes_core_keymem_n2486,
         aes_core_keymem_n2485, aes_core_keymem_n2484, aes_core_keymem_n2483,
         aes_core_keymem_n2482, aes_core_keymem_n2481, aes_core_keymem_n2480,
         aes_core_keymem_n2479, aes_core_keymem_n2478, aes_core_keymem_n2477,
         aes_core_keymem_n2476, aes_core_keymem_n2475, aes_core_keymem_n2474,
         aes_core_keymem_n2473, aes_core_keymem_n2472, aes_core_keymem_n2471,
         aes_core_keymem_n2470, aes_core_keymem_n2469, aes_core_keymem_n2468,
         aes_core_keymem_n2467, aes_core_keymem_n2466, aes_core_keymem_n2465,
         aes_core_keymem_n2464, aes_core_keymem_n2463, aes_core_keymem_n2462,
         aes_core_keymem_n2461, aes_core_keymem_n2460, aes_core_keymem_n2459,
         aes_core_keymem_n2458, aes_core_keymem_n2457, aes_core_keymem_n2456,
         aes_core_keymem_n2455, aes_core_keymem_n2454, aes_core_keymem_n2453,
         aes_core_keymem_n2452, aes_core_keymem_n2451, aes_core_keymem_n2450,
         aes_core_keymem_n2449, aes_core_keymem_n2448, aes_core_keymem_n2447,
         aes_core_keymem_n2446, aes_core_keymem_n2445, aes_core_keymem_n2444,
         aes_core_keymem_n2443, aes_core_keymem_n2442, aes_core_keymem_n2441,
         aes_core_keymem_n2440, aes_core_keymem_n2439, aes_core_keymem_n2438,
         aes_core_keymem_n2437, aes_core_keymem_n2436, aes_core_keymem_n2435,
         aes_core_keymem_n2434, aes_core_keymem_n2433, aes_core_keymem_n2432,
         aes_core_keymem_n2431, aes_core_keymem_n2430, aes_core_keymem_n2429,
         aes_core_keymem_n2428, aes_core_keymem_n2427, aes_core_keymem_n2426,
         aes_core_keymem_n2425, aes_core_keymem_n2424, aes_core_keymem_n2423,
         aes_core_keymem_n2422, aes_core_keymem_n2421, aes_core_keymem_n2420,
         aes_core_keymem_n2419, aes_core_keymem_n2418, aes_core_keymem_n2417,
         aes_core_keymem_n2416, aes_core_keymem_n2415, aes_core_keymem_n2414,
         aes_core_keymem_n2413, aes_core_keymem_n2412, aes_core_keymem_n2411,
         aes_core_keymem_n2410, aes_core_keymem_n2409, aes_core_keymem_n2408,
         aes_core_keymem_n2407, aes_core_keymem_n2406, aes_core_keymem_n2405,
         aes_core_keymem_n2404, aes_core_keymem_n2403, aes_core_keymem_n2402,
         aes_core_keymem_n2401, aes_core_keymem_n2400, aes_core_keymem_n2399,
         aes_core_keymem_n2398, aes_core_keymem_n2397, aes_core_keymem_n2396,
         aes_core_keymem_n2395, aes_core_keymem_n2394, aes_core_keymem_n2393,
         aes_core_keymem_n2392, aes_core_keymem_n2391, aes_core_keymem_n773,
         aes_core_keymem_n770, aes_core_keymem_n767, aes_core_keymem_n764,
         aes_core_keymem_n761, aes_core_keymem_n758, aes_core_keymem_n755,
         aes_core_keymem_n752, aes_core_keymem_n559, aes_core_keymem_n557,
         aes_core_keymem_n554, aes_core_keymem_n544, aes_core_keymem_n30,
         aes_core_keymem_n24, aes_core_keymem_n22, aes_core_keymem_n17,
         aes_core_keymem_n16, aes_core_keymem_n15, aes_core_keymem_n13,
         aes_core_keymem_n12, aes_core_keymem_n11, aes_core_keymem_n10,
         aes_core_keymem_n8, aes_core_keymem_n7, aes_core_keymem_n6,
         aes_core_keymem_n5, aes_core_keymem_n4, aes_core_keymem_n3,
         aes_core_keymem_n2, aes_core_keymem_n1, aes_core_keymem_n2390,
         aes_core_keymem_n2389, aes_core_keymem_n2388, aes_core_keymem_n2387,
         aes_core_keymem_n2386, aes_core_keymem_n2385, aes_core_keymem_n2384,
         aes_core_keymem_n2383, aes_core_keymem_n2382, aes_core_keymem_n2381,
         aes_core_keymem_n2380, aes_core_keymem_n2379, aes_core_keymem_n2378,
         aes_core_keymem_n2377, aes_core_keymem_n2376, aes_core_keymem_n2375,
         aes_core_keymem_n2374, aes_core_keymem_n2373, aes_core_keymem_n2372,
         aes_core_keymem_n2371, aes_core_keymem_n2370, aes_core_keymem_n2369,
         aes_core_keymem_n2368, aes_core_keymem_n2367, aes_core_keymem_n2366,
         aes_core_keymem_n2365, aes_core_keymem_n2364, aes_core_keymem_n2363,
         aes_core_keymem_n2362, aes_core_keymem_n2361, aes_core_keymem_n2360,
         aes_core_keymem_n2359, aes_core_keymem_n2358, aes_core_keymem_n2357,
         aes_core_keymem_n2356, aes_core_keymem_n2355, aes_core_keymem_n2354,
         aes_core_keymem_n2353, aes_core_keymem_n2352, aes_core_keymem_n2351,
         aes_core_keymem_n2350, aes_core_keymem_n2349, aes_core_keymem_n2348,
         aes_core_keymem_n2347, aes_core_keymem_n2346, aes_core_keymem_n2345,
         aes_core_keymem_n2344, aes_core_keymem_n2343, aes_core_keymem_n2342,
         aes_core_keymem_n2341, aes_core_keymem_n2340, aes_core_keymem_n2339,
         aes_core_keymem_n2338, aes_core_keymem_n2337, aes_core_keymem_n2336,
         aes_core_keymem_n2335, aes_core_keymem_n2334, aes_core_keymem_n2333,
         aes_core_keymem_n2332, aes_core_keymem_n2331, aes_core_keymem_n2330,
         aes_core_keymem_n2329, aes_core_keymem_n2328, aes_core_keymem_n2327,
         aes_core_keymem_n2326, aes_core_keymem_n2325, aes_core_keymem_n2324,
         aes_core_keymem_n2323, aes_core_keymem_n2322, aes_core_keymem_n2321,
         aes_core_keymem_n2320, aes_core_keymem_n2319, aes_core_keymem_n2318,
         aes_core_keymem_n2317, aes_core_keymem_n2316, aes_core_keymem_n2315,
         aes_core_keymem_n2314, aes_core_keymem_n2313, aes_core_keymem_n2312,
         aes_core_keymem_n2311, aes_core_keymem_n2310, aes_core_keymem_n2309,
         aes_core_keymem_n2308, aes_core_keymem_n2307, aes_core_keymem_n2306,
         aes_core_keymem_n2305, aes_core_keymem_n2304, aes_core_keymem_n2303,
         aes_core_keymem_n2302, aes_core_keymem_n2301, aes_core_keymem_n2300,
         aes_core_keymem_n2299, aes_core_keymem_n2298, aes_core_keymem_n2297,
         aes_core_keymem_n2296, aes_core_keymem_n2295, aes_core_keymem_n2294,
         aes_core_keymem_n2293, aes_core_keymem_n2292, aes_core_keymem_n2291,
         aes_core_keymem_n2290, aes_core_keymem_n2289, aes_core_keymem_n2288,
         aes_core_keymem_n2287, aes_core_keymem_n2286, aes_core_keymem_n2285,
         aes_core_keymem_n2284, aes_core_keymem_n2283, aes_core_keymem_n2282,
         aes_core_keymem_n2281, aes_core_keymem_n2280, aes_core_keymem_n2279,
         aes_core_keymem_n2278, aes_core_keymem_n2277, aes_core_keymem_n2276,
         aes_core_keymem_n2275, aes_core_keymem_n2274, aes_core_keymem_n2273,
         aes_core_keymem_n2272, aes_core_keymem_n2271, aes_core_keymem_n2270,
         aes_core_keymem_n2269, aes_core_keymem_n2268, aes_core_keymem_n2267,
         aes_core_keymem_n2266, aes_core_keymem_n2265, aes_core_keymem_n2264,
         aes_core_keymem_n2263, aes_core_keymem_n2262, aes_core_keymem_n2261,
         aes_core_keymem_n2260, aes_core_keymem_n2259, aes_core_keymem_n2258,
         aes_core_keymem_n2257, aes_core_keymem_n2256, aes_core_keymem_n2255,
         aes_core_keymem_n2254, aes_core_keymem_n2253, aes_core_keymem_n2252,
         aes_core_keymem_n2251, aes_core_keymem_n2250, aes_core_keymem_n2249,
         aes_core_keymem_n2248, aes_core_keymem_n2247, aes_core_keymem_n2246,
         aes_core_keymem_n2245, aes_core_keymem_n2244, aes_core_keymem_n2243,
         aes_core_keymem_n2242, aes_core_keymem_n2241, aes_core_keymem_n2240,
         aes_core_keymem_n2239, aes_core_keymem_n2238, aes_core_keymem_n2237,
         aes_core_keymem_n2236, aes_core_keymem_n2235, aes_core_keymem_n2234,
         aes_core_keymem_n2233, aes_core_keymem_n2232, aes_core_keymem_n2231,
         aes_core_keymem_n2230, aes_core_keymem_n2229, aes_core_keymem_n2228,
         aes_core_keymem_n2227, aes_core_keymem_n2226, aes_core_keymem_n2225,
         aes_core_keymem_n2224, aes_core_keymem_n2223, aes_core_keymem_n2222,
         aes_core_keymem_n2221, aes_core_keymem_n2220, aes_core_keymem_n2219,
         aes_core_keymem_n2218, aes_core_keymem_n2217, aes_core_keymem_n2216,
         aes_core_keymem_n2215, aes_core_keymem_n2214, aes_core_keymem_n2213,
         aes_core_keymem_n2212, aes_core_keymem_n2211, aes_core_keymem_n2210,
         aes_core_keymem_n2209, aes_core_keymem_n2208, aes_core_keymem_n2207,
         aes_core_keymem_n2206, aes_core_keymem_n2205, aes_core_keymem_n2204,
         aes_core_keymem_n2203, aes_core_keymem_n2202, aes_core_keymem_n2201,
         aes_core_keymem_n2200, aes_core_keymem_n2199, aes_core_keymem_n2198,
         aes_core_keymem_n2197, aes_core_keymem_n2196, aes_core_keymem_n2195,
         aes_core_keymem_n2194, aes_core_keymem_n2193, aes_core_keymem_n2192,
         aes_core_keymem_n2191, aes_core_keymem_n2190, aes_core_keymem_n2189,
         aes_core_keymem_n2188, aes_core_keymem_n2187, aes_core_keymem_n2186,
         aes_core_keymem_n2185, aes_core_keymem_n2184, aes_core_keymem_n2183,
         aes_core_keymem_n2182, aes_core_keymem_n2181, aes_core_keymem_n2180,
         aes_core_keymem_n2179, aes_core_keymem_n2178, aes_core_keymem_n2177,
         aes_core_keymem_n2176, aes_core_keymem_n2175, aes_core_keymem_n2174,
         aes_core_keymem_n2173, aes_core_keymem_n2172, aes_core_keymem_n2171,
         aes_core_keymem_n2170, aes_core_keymem_n2169, aes_core_keymem_n2168,
         aes_core_keymem_n2167, aes_core_keymem_n2166, aes_core_keymem_n2165,
         aes_core_keymem_n2164, aes_core_keymem_n2163, aes_core_keymem_n2162,
         aes_core_keymem_n2161, aes_core_keymem_n2160, aes_core_keymem_n2159,
         aes_core_keymem_n2158, aes_core_keymem_n2157, aes_core_keymem_n2156,
         aes_core_keymem_n2155, aes_core_keymem_n2154, aes_core_keymem_n2153,
         aes_core_keymem_n2152, aes_core_keymem_n2151, aes_core_keymem_n2150,
         aes_core_keymem_n2149, aes_core_keymem_n2148, aes_core_keymem_n2147,
         aes_core_keymem_n2146, aes_core_keymem_n2145, aes_core_keymem_n2144,
         aes_core_keymem_n2143, aes_core_keymem_n2142, aes_core_keymem_n2141,
         aes_core_keymem_n2140, aes_core_keymem_n2139, aes_core_keymem_n2138,
         aes_core_keymem_n2137, aes_core_keymem_n2136, aes_core_keymem_n2135,
         aes_core_keymem_n2134, aes_core_keymem_n2133, aes_core_keymem_n2132,
         aes_core_keymem_n2131, aes_core_keymem_n2130, aes_core_keymem_n2129,
         aes_core_keymem_n2128, aes_core_keymem_n2127, aes_core_keymem_n2126,
         aes_core_keymem_n2125, aes_core_keymem_n2124, aes_core_keymem_n2123,
         aes_core_keymem_n2122, aes_core_keymem_n2121, aes_core_keymem_n2120,
         aes_core_keymem_n2119, aes_core_keymem_n2118, aes_core_keymem_n2117,
         aes_core_keymem_n2116, aes_core_keymem_n2115, aes_core_keymem_n2114,
         aes_core_keymem_n2113, aes_core_keymem_n2112, aes_core_keymem_n2111,
         aes_core_keymem_n2110, aes_core_keymem_n2109, aes_core_keymem_n2108,
         aes_core_keymem_n2107, aes_core_keymem_n2106, aes_core_keymem_n2105,
         aes_core_keymem_n2104, aes_core_keymem_n2103, aes_core_keymem_n2102,
         aes_core_keymem_n2101, aes_core_keymem_n2100, aes_core_keymem_n2099,
         aes_core_keymem_n2098, aes_core_keymem_n2097, aes_core_keymem_n2096,
         aes_core_keymem_n2095, aes_core_keymem_n2094, aes_core_keymem_n2093,
         aes_core_keymem_n2092, aes_core_keymem_n2091, aes_core_keymem_n2090,
         aes_core_keymem_n2089, aes_core_keymem_n2088, aes_core_keymem_n2087,
         aes_core_keymem_n2086, aes_core_keymem_n2085, aes_core_keymem_n2084,
         aes_core_keymem_n2083, aes_core_keymem_n2082, aes_core_keymem_n2081,
         aes_core_keymem_n2080, aes_core_keymem_n2079, aes_core_keymem_n2078,
         aes_core_keymem_n2077, aes_core_keymem_n2076, aes_core_keymem_n2075,
         aes_core_keymem_n2074, aes_core_keymem_n2073, aes_core_keymem_n2072,
         aes_core_keymem_n2071, aes_core_keymem_n2070, aes_core_keymem_n2069,
         aes_core_keymem_n2068, aes_core_keymem_n2067, aes_core_keymem_n2066,
         aes_core_keymem_n2065, aes_core_keymem_n2064, aes_core_keymem_n2063,
         aes_core_keymem_n2062, aes_core_keymem_n2061, aes_core_keymem_n2060,
         aes_core_keymem_n2059, aes_core_keymem_n2058, aes_core_keymem_n2057,
         aes_core_keymem_n2056, aes_core_keymem_n2055, aes_core_keymem_n2054,
         aes_core_keymem_n2053, aes_core_keymem_n2052, aes_core_keymem_n2051,
         aes_core_keymem_n2050, aes_core_keymem_n2049, aes_core_keymem_n2048,
         aes_core_keymem_n2047, aes_core_keymem_n2046, aes_core_keymem_n2045,
         aes_core_keymem_n2044, aes_core_keymem_n2043, aes_core_keymem_n2042,
         aes_core_keymem_n2041, aes_core_keymem_n2040, aes_core_keymem_n2039,
         aes_core_keymem_n2038, aes_core_keymem_n2037, aes_core_keymem_n2036,
         aes_core_keymem_n2035, aes_core_keymem_n2034, aes_core_keymem_n2033,
         aes_core_keymem_n2032, aes_core_keymem_n2031, aes_core_keymem_n2030,
         aes_core_keymem_n2029, aes_core_keymem_n2028, aes_core_keymem_n2027,
         aes_core_keymem_n2026, aes_core_keymem_n2025, aes_core_keymem_n2024,
         aes_core_keymem_n2023, aes_core_keymem_n2022, aes_core_keymem_n2021,
         aes_core_keymem_n2020, aes_core_keymem_n2019, aes_core_keymem_n2018,
         aes_core_keymem_n2017, aes_core_keymem_n2016, aes_core_keymem_n2015,
         aes_core_keymem_n2014, aes_core_keymem_n2013, aes_core_keymem_n2012,
         aes_core_keymem_n2011, aes_core_keymem_n2010, aes_core_keymem_n2009,
         aes_core_keymem_n2008, aes_core_keymem_n2007, aes_core_keymem_n2006,
         aes_core_keymem_n2005, aes_core_keymem_n2004, aes_core_keymem_n2003,
         aes_core_keymem_n2002, aes_core_keymem_n2001, aes_core_keymem_n2000,
         aes_core_keymem_n1999, aes_core_keymem_n1998, aes_core_keymem_n1997,
         aes_core_keymem_n1996, aes_core_keymem_n1995, aes_core_keymem_n1994,
         aes_core_keymem_n1993, aes_core_keymem_n1992, aes_core_keymem_n1991,
         aes_core_keymem_n1990, aes_core_keymem_n1989, aes_core_keymem_n1988,
         aes_core_keymem_n1987, aes_core_keymem_n1986, aes_core_keymem_n1985,
         aes_core_keymem_n1984, aes_core_keymem_n1983, aes_core_keymem_n1982,
         aes_core_keymem_n1981, aes_core_keymem_n1980, aes_core_keymem_n1979,
         aes_core_keymem_n1978, aes_core_keymem_n1977, aes_core_keymem_n1976,
         aes_core_keymem_n1975, aes_core_keymem_n1974, aes_core_keymem_n1973,
         aes_core_keymem_n1972, aes_core_keymem_n1971, aes_core_keymem_n1970,
         aes_core_keymem_n1969, aes_core_keymem_n1968, aes_core_keymem_n1967,
         aes_core_keymem_n1966, aes_core_keymem_n1965, aes_core_keymem_n1964,
         aes_core_keymem_n1963, aes_core_keymem_n1962, aes_core_keymem_n1961,
         aes_core_keymem_n1960, aes_core_keymem_n1959, aes_core_keymem_n1958,
         aes_core_keymem_n1957, aes_core_keymem_n1956, aes_core_keymem_n1955,
         aes_core_keymem_n1954, aes_core_keymem_n1953, aes_core_keymem_n1952,
         aes_core_keymem_n1951, aes_core_keymem_n1950, aes_core_keymem_n1949,
         aes_core_keymem_n1948, aes_core_keymem_n1947, aes_core_keymem_n1946,
         aes_core_keymem_n1945, aes_core_keymem_n1944, aes_core_keymem_n1943,
         aes_core_keymem_n1942, aes_core_keymem_n1941, aes_core_keymem_n1940,
         aes_core_keymem_n1939, aes_core_keymem_n1938, aes_core_keymem_n1937,
         aes_core_keymem_n1936, aes_core_keymem_n1935, aes_core_keymem_n1934,
         aes_core_keymem_n1933, aes_core_keymem_n1932, aes_core_keymem_n1931,
         aes_core_keymem_n1930, aes_core_keymem_n1929, aes_core_keymem_n1928,
         aes_core_keymem_n1927, aes_core_keymem_n1926, aes_core_keymem_n1925,
         aes_core_keymem_n1924, aes_core_keymem_n1923, aes_core_keymem_n1922,
         aes_core_keymem_n1921, aes_core_keymem_n1920, aes_core_keymem_n1919,
         aes_core_keymem_n1918, aes_core_keymem_n1917, aes_core_keymem_n1916,
         aes_core_keymem_n1915, aes_core_keymem_n1914, aes_core_keymem_n1913,
         aes_core_keymem_n1912, aes_core_keymem_n1911, aes_core_keymem_n1910,
         aes_core_keymem_n1909, aes_core_keymem_n1908, aes_core_keymem_n1907,
         aes_core_keymem_n1906, aes_core_keymem_n1905, aes_core_keymem_n1904,
         aes_core_keymem_n1903, aes_core_keymem_n1902, aes_core_keymem_n1901,
         aes_core_keymem_n1900, aes_core_keymem_n1899, aes_core_keymem_n1898,
         aes_core_keymem_n1897, aes_core_keymem_n1896, aes_core_keymem_n1895,
         aes_core_keymem_n1894, aes_core_keymem_n1893, aes_core_keymem_n1892,
         aes_core_keymem_n1891, aes_core_keymem_n1890, aes_core_keymem_n1889,
         aes_core_keymem_n1888, aes_core_keymem_n1887, aes_core_keymem_n1886,
         aes_core_keymem_n1885, aes_core_keymem_n1884, aes_core_keymem_n1883,
         aes_core_keymem_n1882, aes_core_keymem_n1881, aes_core_keymem_n1880,
         aes_core_keymem_n1879, aes_core_keymem_n1878, aes_core_keymem_n1877,
         aes_core_keymem_n1876, aes_core_keymem_n1875, aes_core_keymem_n1874,
         aes_core_keymem_n1873, aes_core_keymem_n1872, aes_core_keymem_n1871,
         aes_core_keymem_n1870, aes_core_keymem_n1869, aes_core_keymem_n1868,
         aes_core_keymem_n1867, aes_core_keymem_n1866, aes_core_keymem_n1865,
         aes_core_keymem_n1864, aes_core_keymem_n1863, aes_core_keymem_n1862,
         aes_core_keymem_n1861, aes_core_keymem_n1860, aes_core_keymem_n1859,
         aes_core_keymem_n1858, aes_core_keymem_n1857, aes_core_keymem_n1856,
         aes_core_keymem_n1855, aes_core_keymem_n1854, aes_core_keymem_n1853,
         aes_core_keymem_n1852, aes_core_keymem_n1851, aes_core_keymem_n1850,
         aes_core_keymem_n1849, aes_core_keymem_n1848, aes_core_keymem_n1847,
         aes_core_keymem_n1846, aes_core_keymem_n1845, aes_core_keymem_n1844,
         aes_core_keymem_n1843, aes_core_keymem_n1842, aes_core_keymem_n1841,
         aes_core_keymem_n1840, aes_core_keymem_n1839, aes_core_keymem_n1838,
         aes_core_keymem_n1837, aes_core_keymem_n1836, aes_core_keymem_n1835,
         aes_core_keymem_n1834, aes_core_keymem_n1833, aes_core_keymem_n1832,
         aes_core_keymem_n1831, aes_core_keymem_n1830, aes_core_keymem_n1829,
         aes_core_keymem_n1828, aes_core_keymem_n1827, aes_core_keymem_n1826,
         aes_core_keymem_n1825, aes_core_keymem_n1824, aes_core_keymem_n1823,
         aes_core_keymem_n1822, aes_core_keymem_n1821, aes_core_keymem_n1820,
         aes_core_keymem_n1819, aes_core_keymem_n1818, aes_core_keymem_n1817,
         aes_core_keymem_n1816, aes_core_keymem_n1815, aes_core_keymem_n1814,
         aes_core_keymem_n1813, aes_core_keymem_n1812, aes_core_keymem_n1811,
         aes_core_keymem_n1810, aes_core_keymem_n1809, aes_core_keymem_n1808,
         aes_core_keymem_n1807, aes_core_keymem_n1806, aes_core_keymem_n1805,
         aes_core_keymem_n1804, aes_core_keymem_n1803, aes_core_keymem_n1802,
         aes_core_keymem_n1801, aes_core_keymem_n1800, aes_core_keymem_n1799,
         aes_core_keymem_n1798, aes_core_keymem_n1797, aes_core_keymem_n1796,
         aes_core_keymem_n1795, aes_core_keymem_n1794, aes_core_keymem_n1793,
         aes_core_keymem_n1792, aes_core_keymem_n1791, aes_core_keymem_n1790,
         aes_core_keymem_n1789, aes_core_keymem_n1788, aes_core_keymem_n1787,
         aes_core_keymem_n1786, aes_core_keymem_n1785, aes_core_keymem_n1784,
         aes_core_keymem_n1783, aes_core_keymem_n1782, aes_core_keymem_n1781,
         aes_core_keymem_n1780, aes_core_keymem_n1779, aes_core_keymem_n1778,
         aes_core_keymem_n1777, aes_core_keymem_n1776, aes_core_keymem_n1775,
         aes_core_keymem_n1774, aes_core_keymem_n1773, aes_core_keymem_n1772,
         aes_core_keymem_n1771, aes_core_keymem_n1770, aes_core_keymem_n1769,
         aes_core_keymem_n1768, aes_core_keymem_n1767, aes_core_keymem_n1766,
         aes_core_keymem_n1765, aes_core_keymem_n1764, aes_core_keymem_n1763,
         aes_core_keymem_n1762, aes_core_keymem_n1761, aes_core_keymem_n1760,
         aes_core_keymem_n1759, aes_core_keymem_n1758, aes_core_keymem_n1757,
         aes_core_keymem_n1756, aes_core_keymem_n1755, aes_core_keymem_n1754,
         aes_core_keymem_n1753, aes_core_keymem_n1752, aes_core_keymem_n1751,
         aes_core_keymem_n1750, aes_core_keymem_n1749, aes_core_keymem_n1748,
         aes_core_keymem_n1747, aes_core_keymem_n1746, aes_core_keymem_n1745,
         aes_core_keymem_n1744, aes_core_keymem_n1743, aes_core_keymem_n1742,
         aes_core_keymem_n1741, aes_core_keymem_n1740, aes_core_keymem_n1739,
         aes_core_keymem_n1738, aes_core_keymem_n1737, aes_core_keymem_n1736,
         aes_core_keymem_n1735, aes_core_keymem_n1734, aes_core_keymem_n1733,
         aes_core_keymem_n1732, aes_core_keymem_n1731, aes_core_keymem_n1730,
         aes_core_keymem_n1729, aes_core_keymem_n1728, aes_core_keymem_n1727,
         aes_core_keymem_n1726, aes_core_keymem_n1725, aes_core_keymem_n1724,
         aes_core_keymem_n1723, aes_core_keymem_n1722, aes_core_keymem_n1721,
         aes_core_keymem_n1720, aes_core_keymem_n1719, aes_core_keymem_n1718,
         aes_core_keymem_n1717, aes_core_keymem_n1716, aes_core_keymem_n1715,
         aes_core_keymem_n1714, aes_core_keymem_n1713, aes_core_keymem_n1712,
         aes_core_keymem_n1711, aes_core_keymem_n1710, aes_core_keymem_n1709,
         aes_core_keymem_n1708, aes_core_keymem_n1707, aes_core_keymem_n1706,
         aes_core_keymem_n1705, aes_core_keymem_n1704, aes_core_keymem_n1703,
         aes_core_keymem_n1702, aes_core_keymem_n1701, aes_core_keymem_n1700,
         aes_core_keymem_n1699, aes_core_keymem_n1698, aes_core_keymem_n1697,
         aes_core_keymem_n1696, aes_core_keymem_n1695, aes_core_keymem_n1694,
         aes_core_keymem_n1693, aes_core_keymem_n1692, aes_core_keymem_n1691,
         aes_core_keymem_n1690, aes_core_keymem_n1689, aes_core_keymem_n1688,
         aes_core_keymem_n1687, aes_core_keymem_n1686, aes_core_keymem_n1685,
         aes_core_keymem_n1684, aes_core_keymem_n1683, aes_core_keymem_n1682,
         aes_core_keymem_n1681, aes_core_keymem_n1680, aes_core_keymem_n1679,
         aes_core_keymem_n1678, aes_core_keymem_n1677, aes_core_keymem_n1676,
         aes_core_keymem_n1675, aes_core_keymem_n1674, aes_core_keymem_n1673,
         aes_core_keymem_n1672, aes_core_keymem_n1671, aes_core_keymem_n1670,
         aes_core_keymem_n1669, aes_core_keymem_n1668, aes_core_keymem_n1667,
         aes_core_keymem_n1666, aes_core_keymem_n1665, aes_core_keymem_n1664,
         aes_core_keymem_n1663, aes_core_keymem_n1662, aes_core_keymem_n1661,
         aes_core_keymem_n1660, aes_core_keymem_n1659, aes_core_keymem_n1658,
         aes_core_keymem_n1657, aes_core_keymem_n1656, aes_core_keymem_n1655,
         aes_core_keymem_n1654, aes_core_keymem_n1653, aes_core_keymem_n1652,
         aes_core_keymem_n1651, aes_core_keymem_n1650, aes_core_keymem_n1649,
         aes_core_keymem_n1648, aes_core_keymem_n1647, aes_core_keymem_n1646,
         aes_core_keymem_n1645, aes_core_keymem_n1644, aes_core_keymem_n1643,
         aes_core_keymem_n1642, aes_core_keymem_n1641, aes_core_keymem_n1640,
         aes_core_keymem_n1639, aes_core_keymem_n1638, aes_core_keymem_n1637,
         aes_core_keymem_n1636, aes_core_keymem_n1635, aes_core_keymem_n1634,
         aes_core_keymem_n1633, aes_core_keymem_n1632, aes_core_keymem_n1631,
         aes_core_keymem_n1630, aes_core_keymem_n1629, aes_core_keymem_n1628,
         aes_core_keymem_n1627, aes_core_keymem_n1626, aes_core_keymem_n1625,
         aes_core_keymem_n1624, aes_core_keymem_n1623, aes_core_keymem_n1622,
         aes_core_keymem_n1621, aes_core_keymem_n1620, aes_core_keymem_n1619,
         aes_core_keymem_n1618, aes_core_keymem_n1617, aes_core_keymem_n1616,
         aes_core_keymem_n1615, aes_core_keymem_n1614, aes_core_keymem_n1613,
         aes_core_keymem_n1612, aes_core_keymem_n1611, aes_core_keymem_n1610,
         aes_core_keymem_n1609, aes_core_keymem_n1608, aes_core_keymem_n1607,
         aes_core_keymem_n1606, aes_core_keymem_n1605, aes_core_keymem_n1604,
         aes_core_keymem_n1603, aes_core_keymem_n1602, aes_core_keymem_n1601,
         aes_core_keymem_n1600, aes_core_keymem_n1599, aes_core_keymem_n1598,
         aes_core_keymem_n1597, aes_core_keymem_n1596, aes_core_keymem_n1595,
         aes_core_keymem_n1594, aes_core_keymem_n1593, aes_core_keymem_n1592,
         aes_core_keymem_n1591, aes_core_keymem_n1590, aes_core_keymem_n1589,
         aes_core_keymem_n1588, aes_core_keymem_n1587, aes_core_keymem_n1586,
         aes_core_keymem_n1585, aes_core_keymem_n1584, aes_core_keymem_n1583,
         aes_core_keymem_n1582, aes_core_keymem_n1581, aes_core_keymem_n1580,
         aes_core_keymem_n1579, aes_core_keymem_n1578, aes_core_keymem_n1577,
         aes_core_keymem_n1576, aes_core_keymem_n1575, aes_core_keymem_n1574,
         aes_core_keymem_n1573, aes_core_keymem_n1572, aes_core_keymem_n1571,
         aes_core_keymem_n1570, aes_core_keymem_n1569, aes_core_keymem_n1568,
         aes_core_keymem_n1567, aes_core_keymem_n1566, aes_core_keymem_n1565,
         aes_core_keymem_n1564, aes_core_keymem_n1563, aes_core_keymem_n1562,
         aes_core_keymem_n1561, aes_core_keymem_n1560, aes_core_keymem_n1559,
         aes_core_keymem_n1558, aes_core_keymem_n1557, aes_core_keymem_n1556,
         aes_core_keymem_n1555, aes_core_keymem_n1554, aes_core_keymem_n1553,
         aes_core_keymem_n1552, aes_core_keymem_n1551, aes_core_keymem_n1550,
         aes_core_keymem_n1549, aes_core_keymem_n1548, aes_core_keymem_n1547,
         aes_core_keymem_n1546, aes_core_keymem_n1545, aes_core_keymem_n1544,
         aes_core_keymem_n1543, aes_core_keymem_n1542, aes_core_keymem_n1541,
         aes_core_keymem_n1540, aes_core_keymem_n1539, aes_core_keymem_n1538,
         aes_core_keymem_n1537, aes_core_keymem_n1536, aes_core_keymem_n1535,
         aes_core_keymem_n1534, aes_core_keymem_n1533, aes_core_keymem_n1532,
         aes_core_keymem_n1531, aes_core_keymem_n1530, aes_core_keymem_n1529,
         aes_core_keymem_n1528, aes_core_keymem_n1527, aes_core_keymem_n1526,
         aes_core_keymem_n1525, aes_core_keymem_n1524, aes_core_keymem_n1523,
         aes_core_keymem_n1522, aes_core_keymem_n1521, aes_core_keymem_n1520,
         aes_core_keymem_n1519, aes_core_keymem_n1518, aes_core_keymem_n1517,
         aes_core_keymem_n1516, aes_core_keymem_n1515, aes_core_keymem_n1514,
         aes_core_keymem_n1513, aes_core_keymem_n1512, aes_core_keymem_n1511,
         aes_core_keymem_n1510, aes_core_keymem_n1509, aes_core_keymem_n1508,
         aes_core_keymem_n1507, aes_core_keymem_n1506, aes_core_keymem_n1505,
         aes_core_keymem_n1504, aes_core_keymem_n1503, aes_core_keymem_n1502,
         aes_core_keymem_n1501, aes_core_keymem_n1500, aes_core_keymem_n1499,
         aes_core_keymem_n1498, aes_core_keymem_n1497, aes_core_keymem_n1496,
         aes_core_keymem_n1495, aes_core_keymem_n1494, aes_core_keymem_n1493,
         aes_core_keymem_n1492, aes_core_keymem_n1491, aes_core_keymem_n1490,
         aes_core_keymem_n1489, aes_core_keymem_n1488, aes_core_keymem_n1487,
         aes_core_keymem_n1486, aes_core_keymem_n1485, aes_core_keymem_n1484,
         aes_core_keymem_n1483, aes_core_keymem_n1482, aes_core_keymem_n1481,
         aes_core_keymem_n1480, aes_core_keymem_n1479, aes_core_keymem_n1478,
         aes_core_keymem_n1477, aes_core_keymem_n1476, aes_core_keymem_n1475,
         aes_core_keymem_n1474, aes_core_keymem_n1473, aes_core_keymem_n1472,
         aes_core_keymem_n1471, aes_core_keymem_n1470, aes_core_keymem_n1469,
         aes_core_keymem_n1468, aes_core_keymem_n1467, aes_core_keymem_n1466,
         aes_core_keymem_n1465, aes_core_keymem_n1464, aes_core_keymem_n1463,
         aes_core_keymem_n1462, aes_core_keymem_n1461, aes_core_keymem_n1460,
         aes_core_keymem_n1459, aes_core_keymem_n1458, aes_core_keymem_n1457,
         aes_core_keymem_n1456, aes_core_keymem_n1455, aes_core_keymem_n1454,
         aes_core_keymem_n1453, aes_core_keymem_n1452, aes_core_keymem_n1451,
         aes_core_keymem_n1450, aes_core_keymem_n1449, aes_core_keymem_n1448,
         aes_core_keymem_n1447, aes_core_keymem_n1446, aes_core_keymem_n1445,
         aes_core_keymem_n1444, aes_core_keymem_n1443, aes_core_keymem_n1442,
         aes_core_keymem_n1441, aes_core_keymem_n1440, aes_core_keymem_n1439,
         aes_core_keymem_n1438, aes_core_keymem_n1437, aes_core_keymem_n1436,
         aes_core_keymem_n1435, aes_core_keymem_n1434, aes_core_keymem_n1433,
         aes_core_keymem_n1432, aes_core_keymem_n1431, aes_core_keymem_n1430,
         aes_core_keymem_n1429, aes_core_keymem_n1428, aes_core_keymem_n1427,
         aes_core_keymem_n1426, aes_core_keymem_n1425, aes_core_keymem_n1424,
         aes_core_keymem_n1423, aes_core_keymem_n1422, aes_core_keymem_n1421,
         aes_core_keymem_n1420, aes_core_keymem_n1419, aes_core_keymem_n1418,
         aes_core_keymem_n1417, aes_core_keymem_n1416, aes_core_keymem_n1415,
         aes_core_keymem_n1414, aes_core_keymem_n1413, aes_core_keymem_n1412,
         aes_core_keymem_n1411, aes_core_keymem_n1410, aes_core_keymem_n1409,
         aes_core_keymem_n1408, aes_core_keymem_n1407, aes_core_keymem_n1406,
         aes_core_keymem_n1405, aes_core_keymem_n1404, aes_core_keymem_n1403,
         aes_core_keymem_n1402, aes_core_keymem_n1401, aes_core_keymem_n1400,
         aes_core_keymem_n1399, aes_core_keymem_n1398, aes_core_keymem_n1397,
         aes_core_keymem_n1396, aes_core_keymem_n1395, aes_core_keymem_n1394,
         aes_core_keymem_n1393, aes_core_keymem_n1392, aes_core_keymem_n1391,
         aes_core_keymem_n1390, aes_core_keymem_n1389, aes_core_keymem_n1388,
         aes_core_keymem_n1387, aes_core_keymem_n1386, aes_core_keymem_n1385,
         aes_core_keymem_n1384, aes_core_keymem_n1383, aes_core_keymem_n1382,
         aes_core_keymem_n1381, aes_core_keymem_n1380, aes_core_keymem_n1379,
         aes_core_keymem_n1378, aes_core_keymem_n1377, aes_core_keymem_n1376,
         aes_core_keymem_n1375, aes_core_keymem_n1374, aes_core_keymem_n1373,
         aes_core_keymem_n1372, aes_core_keymem_n1371, aes_core_keymem_n1370,
         aes_core_keymem_n1369, aes_core_keymem_n1368, aes_core_keymem_n1367,
         aes_core_keymem_n1366, aes_core_keymem_n1365, aes_core_keymem_n1364,
         aes_core_keymem_n1363, aes_core_keymem_n1362, aes_core_keymem_n1361,
         aes_core_keymem_n1360, aes_core_keymem_n1359, aes_core_keymem_n1358,
         aes_core_keymem_n1357, aes_core_keymem_n1356, aes_core_keymem_n1355,
         aes_core_keymem_n1354, aes_core_keymem_n1353, aes_core_keymem_n1352,
         aes_core_keymem_n1351, aes_core_keymem_n1350, aes_core_keymem_n1349,
         aes_core_keymem_n1348, aes_core_keymem_n1347, aes_core_keymem_n1346,
         aes_core_keymem_n1345, aes_core_keymem_n1344, aes_core_keymem_n1343,
         aes_core_keymem_n1342, aes_core_keymem_n1341, aes_core_keymem_n1340,
         aes_core_keymem_n1339, aes_core_keymem_n1338, aes_core_keymem_n1337,
         aes_core_keymem_n1336, aes_core_keymem_n1335, aes_core_keymem_n1334,
         aes_core_keymem_n1333, aes_core_keymem_n1332, aes_core_keymem_n1331,
         aes_core_keymem_n1330, aes_core_keymem_n1329, aes_core_keymem_n1328,
         aes_core_keymem_n1327, aes_core_keymem_n1326, aes_core_keymem_n1325,
         aes_core_keymem_n1324, aes_core_keymem_n1323, aes_core_keymem_n1322,
         aes_core_keymem_n1321, aes_core_keymem_n1320, aes_core_keymem_n1319,
         aes_core_keymem_n1318, aes_core_keymem_n1317, aes_core_keymem_n1316,
         aes_core_keymem_n1315, aes_core_keymem_n1314, aes_core_keymem_n1313,
         aes_core_keymem_n1312, aes_core_keymem_n1311, aes_core_keymem_n1310,
         aes_core_keymem_n1309, aes_core_keymem_n1308, aes_core_keymem_n1307,
         aes_core_keymem_n1306, aes_core_keymem_n1305, aes_core_keymem_n1304,
         aes_core_keymem_n1303, aes_core_keymem_n1302, aes_core_keymem_n1301,
         aes_core_keymem_n1300, aes_core_keymem_n1299, aes_core_keymem_n1298,
         aes_core_keymem_n1297, aes_core_keymem_n1296, aes_core_keymem_n1295,
         aes_core_keymem_n1294, aes_core_keymem_n1293, aes_core_keymem_n1292,
         aes_core_keymem_n1291, aes_core_keymem_n1290, aes_core_keymem_n1289,
         aes_core_keymem_n1288, aes_core_keymem_n1287, aes_core_keymem_n1286,
         aes_core_keymem_n1285, aes_core_keymem_n1284, aes_core_keymem_n1283,
         aes_core_keymem_n1282, aes_core_keymem_n1281, aes_core_keymem_n1280,
         aes_core_keymem_n1279, aes_core_keymem_n1278, aes_core_keymem_n1277,
         aes_core_keymem_n1276, aes_core_keymem_n1275, aes_core_keymem_n1274,
         aes_core_keymem_n1273, aes_core_keymem_n1272, aes_core_keymem_n1271,
         aes_core_keymem_n1270, aes_core_keymem_n1269, aes_core_keymem_n1268,
         aes_core_keymem_n1267, aes_core_keymem_n1266, aes_core_keymem_n1265,
         aes_core_keymem_n1264, aes_core_keymem_n1263, aes_core_keymem_n1262,
         aes_core_keymem_n1261, aes_core_keymem_n1260, aes_core_keymem_n1259,
         aes_core_keymem_n1258, aes_core_keymem_n1257, aes_core_keymem_n1256,
         aes_core_keymem_n1255, aes_core_keymem_n1254, aes_core_keymem_n1253,
         aes_core_keymem_n1252, aes_core_keymem_n1251, aes_core_keymem_n1250,
         aes_core_keymem_n1249, aes_core_keymem_n1248, aes_core_keymem_n1247,
         aes_core_keymem_n1246, aes_core_keymem_n1245, aes_core_keymem_n1244,
         aes_core_keymem_n1243, aes_core_keymem_n1242, aes_core_keymem_n1241,
         aes_core_keymem_n1240, aes_core_keymem_n1239, aes_core_keymem_n1238,
         aes_core_keymem_n1237, aes_core_keymem_n1236, aes_core_keymem_n1235,
         aes_core_keymem_n1234, aes_core_keymem_n1233, aes_core_keymem_n1232,
         aes_core_keymem_n1231, aes_core_keymem_n1230, aes_core_keymem_n1229,
         aes_core_keymem_n1228, aes_core_keymem_n1227, aes_core_keymem_n1226,
         aes_core_keymem_n1225, aes_core_keymem_n1224, aes_core_keymem_n1223,
         aes_core_keymem_n1222, aes_core_keymem_n1221, aes_core_keymem_n1220,
         aes_core_keymem_n1219, aes_core_keymem_n1218, aes_core_keymem_n1217,
         aes_core_keymem_n1216, aes_core_keymem_n1215, aes_core_keymem_n1214,
         aes_core_keymem_n1213, aes_core_keymem_n1212, aes_core_keymem_n1211,
         aes_core_keymem_n1210, aes_core_keymem_n1209, aes_core_keymem_n1208,
         aes_core_keymem_n1207, aes_core_keymem_n1206, aes_core_keymem_n1205,
         aes_core_keymem_n1204, aes_core_keymem_n1203, aes_core_keymem_n1202,
         aes_core_keymem_n1201, aes_core_keymem_n1200, aes_core_keymem_n1199,
         aes_core_keymem_n1198, aes_core_keymem_n1197, aes_core_keymem_n1196,
         aes_core_keymem_n1195, aes_core_keymem_n1194, aes_core_keymem_n1193,
         aes_core_keymem_n1192, aes_core_keymem_n1191, aes_core_keymem_n1190,
         aes_core_keymem_n1189, aes_core_keymem_n1188, aes_core_keymem_n1187,
         aes_core_keymem_n1186, aes_core_keymem_n1185, aes_core_keymem_n1184,
         aes_core_keymem_n1183, aes_core_keymem_n1182, aes_core_keymem_n1181,
         aes_core_keymem_n1180, aes_core_keymem_n1179, aes_core_keymem_n1178,
         aes_core_keymem_n1177, aes_core_keymem_n1176, aes_core_keymem_n1175,
         aes_core_keymem_n1174, aes_core_keymem_n1173, aes_core_keymem_n1172,
         aes_core_keymem_n1171, aes_core_keymem_n1170, aes_core_keymem_n1169,
         aes_core_keymem_n1168, aes_core_keymem_n1167, aes_core_keymem_n1166,
         aes_core_keymem_n1165, aes_core_keymem_n1164, aes_core_keymem_n1163,
         aes_core_keymem_n1162, aes_core_keymem_n1161, aes_core_keymem_n1160,
         aes_core_keymem_n1159, aes_core_keymem_n1158, aes_core_keymem_n1157,
         aes_core_keymem_n1156, aes_core_keymem_n1155, aes_core_keymem_n1154,
         aes_core_keymem_n1153, aes_core_keymem_n1152, aes_core_keymem_n1151,
         aes_core_keymem_n1150, aes_core_keymem_n1149, aes_core_keymem_n1148,
         aes_core_keymem_n1147, aes_core_keymem_n1146, aes_core_keymem_n1145,
         aes_core_keymem_n1144, aes_core_keymem_n1143, aes_core_keymem_n1142,
         aes_core_keymem_n1141, aes_core_keymem_n1140, aes_core_keymem_n1139,
         aes_core_keymem_n1138, aes_core_keymem_n1137, aes_core_keymem_n1136,
         aes_core_keymem_n1135, aes_core_keymem_n1134, aes_core_keymem_n1133,
         aes_core_keymem_n1132, aes_core_keymem_n1131, aes_core_keymem_n1130,
         aes_core_keymem_n1129, aes_core_keymem_n1128, aes_core_keymem_n1127,
         aes_core_keymem_n1126, aes_core_keymem_n1125, aes_core_keymem_n1124,
         aes_core_keymem_n1123, aes_core_keymem_n1122, aes_core_keymem_n1121,
         aes_core_keymem_n1120, aes_core_keymem_n1119, aes_core_keymem_n1118,
         aes_core_keymem_n1117, aes_core_keymem_n1116, aes_core_keymem_n1115,
         aes_core_keymem_n1114, aes_core_keymem_n1113, aes_core_keymem_n1112,
         aes_core_keymem_n1111, aes_core_keymem_n1110, aes_core_keymem_n1109,
         aes_core_keymem_n1108, aes_core_keymem_n1107, aes_core_keymem_n1106,
         aes_core_keymem_n1105, aes_core_keymem_n1104, aes_core_keymem_n1103,
         aes_core_keymem_n1102, aes_core_keymem_n1101, aes_core_keymem_n1100,
         aes_core_keymem_n1099, aes_core_keymem_n1098, aes_core_keymem_n1097,
         aes_core_keymem_n1096, aes_core_keymem_n1095, aes_core_keymem_n1094,
         aes_core_keymem_n1093, aes_core_keymem_n1092, aes_core_keymem_n1091,
         aes_core_keymem_n1090, aes_core_keymem_n1089, aes_core_keymem_n1088,
         aes_core_keymem_n1087, aes_core_keymem_n1086, aes_core_keymem_n1085,
         aes_core_keymem_n1084, aes_core_keymem_n1083, aes_core_keymem_n1082,
         aes_core_keymem_n1081, aes_core_keymem_n1080, aes_core_keymem_n1079,
         aes_core_keymem_n1078, aes_core_keymem_n1077, aes_core_keymem_n1076,
         aes_core_keymem_n1075, aes_core_keymem_n1074, aes_core_keymem_n1073,
         aes_core_keymem_n1072, aes_core_keymem_n1071, aes_core_keymem_n1070,
         aes_core_keymem_n1069, aes_core_keymem_n1068, aes_core_keymem_n1067,
         aes_core_keymem_n1066, aes_core_keymem_n1065, aes_core_keymem_n1064,
         aes_core_keymem_n1063, aes_core_keymem_n1062, aes_core_keymem_n1061,
         aes_core_keymem_n1060, aes_core_keymem_n1059, aes_core_keymem_n1058,
         aes_core_keymem_n1057, aes_core_keymem_n1056, aes_core_keymem_n1055,
         aes_core_keymem_n1054, aes_core_keymem_n1053, aes_core_keymem_n1052,
         aes_core_keymem_n1051, aes_core_keymem_n1050, aes_core_keymem_n1049,
         aes_core_keymem_n1048, aes_core_keymem_n1047, aes_core_keymem_n1046,
         aes_core_keymem_n1045, aes_core_keymem_n1044, aes_core_keymem_n1043,
         aes_core_keymem_n1042, aes_core_keymem_n1041, aes_core_keymem_n1040,
         aes_core_keymem_n1039, aes_core_keymem_n1038, aes_core_keymem_n1037,
         aes_core_keymem_n1036, aes_core_keymem_n1035, aes_core_keymem_n1034,
         aes_core_keymem_n1033, aes_core_keymem_n1032, aes_core_keymem_n1031,
         aes_core_keymem_n1030, aes_core_keymem_n1029, aes_core_keymem_n1028,
         aes_core_keymem_n1027, aes_core_keymem_n1026, aes_core_keymem_n1025,
         aes_core_keymem_n1024, aes_core_keymem_n1023, aes_core_keymem_n1022,
         aes_core_keymem_n1021, aes_core_keymem_n1020, aes_core_keymem_n1019,
         aes_core_keymem_n1018, aes_core_keymem_n1017, aes_core_keymem_n1016,
         aes_core_keymem_n1015, aes_core_keymem_n1014, aes_core_keymem_n1013,
         aes_core_keymem_n1012, aes_core_keymem_n1011, aes_core_keymem_n1010,
         aes_core_keymem_n1009, aes_core_keymem_n1008, aes_core_keymem_n1007,
         aes_core_keymem_n1006, aes_core_keymem_n1005, aes_core_keymem_n1004,
         aes_core_keymem_n1003, aes_core_keymem_n1002, aes_core_keymem_n1001,
         aes_core_keymem_n1000, aes_core_keymem_n999, aes_core_keymem_n998,
         aes_core_keymem_n997, aes_core_keymem_n996, aes_core_keymem_n995,
         aes_core_keymem_n994, aes_core_keymem_n993, aes_core_keymem_n992,
         aes_core_keymem_n991, aes_core_keymem_n990, aes_core_keymem_n989,
         aes_core_keymem_n988, aes_core_keymem_n987, aes_core_keymem_n986,
         aes_core_keymem_n985, aes_core_keymem_n984, aes_core_keymem_n983,
         aes_core_keymem_n982, aes_core_keymem_n981, aes_core_keymem_n980,
         aes_core_keymem_n979, aes_core_keymem_n978, aes_core_keymem_n977,
         aes_core_keymem_n976, aes_core_keymem_n975, aes_core_keymem_n974,
         aes_core_keymem_n973, aes_core_keymem_n972, aes_core_keymem_n971,
         aes_core_keymem_n970, aes_core_keymem_n969, aes_core_keymem_n968,
         aes_core_keymem_n967, aes_core_keymem_n966, aes_core_keymem_n965,
         aes_core_keymem_n964, aes_core_keymem_n963, aes_core_keymem_n962,
         aes_core_keymem_n961, aes_core_keymem_n960, aes_core_keymem_n959,
         aes_core_keymem_n958, aes_core_keymem_n957, aes_core_keymem_n956,
         aes_core_keymem_n955, aes_core_keymem_n954, aes_core_keymem_n953,
         aes_core_keymem_n952, aes_core_keymem_n951, aes_core_keymem_n950,
         aes_core_keymem_n949, aes_core_keymem_n948, aes_core_keymem_n947,
         aes_core_keymem_n946, aes_core_keymem_n945, aes_core_keymem_n944,
         aes_core_keymem_n943, aes_core_keymem_n942, aes_core_keymem_n941,
         aes_core_keymem_n940, aes_core_keymem_n939, aes_core_keymem_n938,
         aes_core_keymem_n937, aes_core_keymem_n936, aes_core_keymem_n935,
         aes_core_keymem_n934, aes_core_keymem_n933, aes_core_keymem_n932,
         aes_core_keymem_n931, aes_core_keymem_n930, aes_core_keymem_n929,
         aes_core_keymem_n928, aes_core_keymem_n927, aes_core_keymem_n926,
         aes_core_keymem_n925, aes_core_keymem_n924, aes_core_keymem_n923,
         aes_core_keymem_n922, aes_core_keymem_n921, aes_core_keymem_n920,
         aes_core_keymem_n919, aes_core_keymem_n918, aes_core_keymem_n917,
         aes_core_keymem_n916, aes_core_keymem_n915, aes_core_keymem_n914,
         aes_core_keymem_n913, aes_core_keymem_n912, aes_core_keymem_n911,
         aes_core_keymem_n910, aes_core_keymem_n909, aes_core_keymem_n908,
         aes_core_keymem_n907, aes_core_keymem_n906, aes_core_keymem_n905,
         aes_core_keymem_n904, aes_core_keymem_n903, aes_core_keymem_n902,
         aes_core_keymem_n901, aes_core_keymem_n900, aes_core_keymem_n899,
         aes_core_keymem_n898, aes_core_keymem_n897, aes_core_keymem_n896,
         aes_core_keymem_n895, aes_core_keymem_n894, aes_core_keymem_n893,
         aes_core_keymem_n892, aes_core_keymem_n891, aes_core_keymem_n890,
         aes_core_keymem_n889, aes_core_keymem_n888, aes_core_keymem_n887,
         aes_core_keymem_n886, aes_core_keymem_n885, aes_core_keymem_n884,
         aes_core_keymem_n883, aes_core_keymem_n882, aes_core_keymem_n881,
         aes_core_keymem_n880, aes_core_keymem_n879, aes_core_keymem_n878,
         aes_core_keymem_n877, aes_core_keymem_n876, aes_core_keymem_n875,
         aes_core_keymem_n874, aes_core_keymem_n873, aes_core_keymem_n872,
         aes_core_keymem_n871, aes_core_keymem_n870, aes_core_keymem_n869,
         aes_core_keymem_n868, aes_core_keymem_n867, aes_core_keymem_n866,
         aes_core_keymem_n865, aes_core_keymem_n864, aes_core_keymem_n863,
         aes_core_keymem_n862, aes_core_keymem_n861, aes_core_keymem_n860,
         aes_core_keymem_n859, aes_core_keymem_n858, aes_core_keymem_n857,
         aes_core_keymem_n856, aes_core_keymem_n855, aes_core_keymem_n854,
         aes_core_keymem_n853, aes_core_keymem_n852, aes_core_keymem_n851,
         aes_core_keymem_n850, aes_core_keymem_n849, aes_core_keymem_n848,
         aes_core_keymem_n847, aes_core_keymem_n846, aes_core_keymem_n845,
         aes_core_keymem_n844, aes_core_keymem_n843, aes_core_keymem_n842,
         aes_core_keymem_n841, aes_core_keymem_n840, aes_core_keymem_n839,
         aes_core_keymem_n838, aes_core_keymem_n837, aes_core_keymem_n836,
         aes_core_keymem_n835, aes_core_keymem_n834, aes_core_keymem_n833,
         aes_core_keymem_n832, aes_core_keymem_n831, aes_core_keymem_n830,
         aes_core_keymem_n829, aes_core_keymem_n828, aes_core_keymem_n827,
         aes_core_keymem_n826, aes_core_keymem_n825, aes_core_keymem_n824,
         aes_core_keymem_n823, aes_core_keymem_n822, aes_core_keymem_n821,
         aes_core_keymem_n820, aes_core_keymem_n819, aes_core_keymem_n818,
         aes_core_keymem_n817, aes_core_keymem_n816, aes_core_keymem_n815,
         aes_core_keymem_n814, aes_core_keymem_n813, aes_core_keymem_n812,
         aes_core_keymem_n811, aes_core_keymem_n810, aes_core_keymem_n809,
         aes_core_keymem_n808, aes_core_keymem_n807, aes_core_keymem_n806,
         aes_core_keymem_n805, aes_core_keymem_n804, aes_core_keymem_n803,
         aes_core_keymem_n802, aes_core_keymem_n801, aes_core_keymem_n800,
         aes_core_keymem_n799, aes_core_keymem_n798, aes_core_keymem_n797,
         aes_core_keymem_n796, aes_core_keymem_n795, aes_core_keymem_n794,
         aes_core_keymem_n793, aes_core_keymem_n792, aes_core_keymem_n791,
         aes_core_keymem_n790, aes_core_keymem_n789, aes_core_keymem_n788,
         aes_core_keymem_n787, aes_core_keymem_n786, aes_core_keymem_n785,
         aes_core_keymem_n784, aes_core_keymem_n783, aes_core_keymem_n782,
         aes_core_keymem_n781, aes_core_keymem_n780, aes_core_keymem_n779,
         aes_core_keymem_n778, aes_core_keymem_n777, aes_core_keymem_n776,
         aes_core_keymem_n775, aes_core_keymem_n774, aes_core_keymem_n772,
         aes_core_keymem_n771, aes_core_keymem_n769, aes_core_keymem_n768,
         aes_core_keymem_n766, aes_core_keymem_n765, aes_core_keymem_n763,
         aes_core_keymem_n762, aes_core_keymem_n760, aes_core_keymem_n759,
         aes_core_keymem_n757, aes_core_keymem_n756, aes_core_keymem_n754,
         aes_core_keymem_n753, aes_core_keymem_n751, aes_core_keymem_n750,
         aes_core_keymem_n749, aes_core_keymem_n748, aes_core_keymem_n747,
         aes_core_keymem_n746, aes_core_keymem_n745, aes_core_keymem_n744,
         aes_core_keymem_n743, aes_core_keymem_n742, aes_core_keymem_n741,
         aes_core_keymem_n740, aes_core_keymem_n739, aes_core_keymem_n738,
         aes_core_keymem_n737, aes_core_keymem_n736, aes_core_keymem_n735,
         aes_core_keymem_n734, aes_core_keymem_n733, aes_core_keymem_n732,
         aes_core_keymem_n731, aes_core_keymem_n730, aes_core_keymem_n729,
         aes_core_keymem_n728, aes_core_keymem_n727, aes_core_keymem_n726,
         aes_core_keymem_n725, aes_core_keymem_n724, aes_core_keymem_n723,
         aes_core_keymem_n722, aes_core_keymem_n721, aes_core_keymem_n720,
         aes_core_keymem_n719, aes_core_keymem_n718, aes_core_keymem_n717,
         aes_core_keymem_n716, aes_core_keymem_n715, aes_core_keymem_n714,
         aes_core_keymem_n713, aes_core_keymem_n712, aes_core_keymem_n711,
         aes_core_keymem_n710, aes_core_keymem_n709, aes_core_keymem_n708,
         aes_core_keymem_n707, aes_core_keymem_n706, aes_core_keymem_n705,
         aes_core_keymem_n704, aes_core_keymem_n703, aes_core_keymem_n702,
         aes_core_keymem_n701, aes_core_keymem_n700, aes_core_keymem_n699,
         aes_core_keymem_n698, aes_core_keymem_n697, aes_core_keymem_n696,
         aes_core_keymem_n695, aes_core_keymem_n694, aes_core_keymem_n693,
         aes_core_keymem_n692, aes_core_keymem_n691, aes_core_keymem_n690,
         aes_core_keymem_n689, aes_core_keymem_n688, aes_core_keymem_n687,
         aes_core_keymem_n686, aes_core_keymem_n685, aes_core_keymem_n684,
         aes_core_keymem_n683, aes_core_keymem_n682, aes_core_keymem_n681,
         aes_core_keymem_n680, aes_core_keymem_n679, aes_core_keymem_n678,
         aes_core_keymem_n677, aes_core_keymem_n676, aes_core_keymem_n675,
         aes_core_keymem_n674, aes_core_keymem_n673, aes_core_keymem_n672,
         aes_core_keymem_n671, aes_core_keymem_n670, aes_core_keymem_n669,
         aes_core_keymem_n668, aes_core_keymem_n667, aes_core_keymem_n666,
         aes_core_keymem_n665, aes_core_keymem_n664, aes_core_keymem_n663,
         aes_core_keymem_n662, aes_core_keymem_n661, aes_core_keymem_n660,
         aes_core_keymem_n659, aes_core_keymem_n658, aes_core_keymem_n657,
         aes_core_keymem_n656, aes_core_keymem_n655, aes_core_keymem_n654,
         aes_core_keymem_n653, aes_core_keymem_n652, aes_core_keymem_n651,
         aes_core_keymem_n650, aes_core_keymem_n649, aes_core_keymem_n648,
         aes_core_keymem_n647, aes_core_keymem_n646, aes_core_keymem_n645,
         aes_core_keymem_n644, aes_core_keymem_n643, aes_core_keymem_n642,
         aes_core_keymem_n641, aes_core_keymem_n640, aes_core_keymem_n639,
         aes_core_keymem_n638, aes_core_keymem_n637, aes_core_keymem_n636,
         aes_core_keymem_n635, aes_core_keymem_n634, aes_core_keymem_n633,
         aes_core_keymem_n632, aes_core_keymem_n631, aes_core_keymem_n630,
         aes_core_keymem_n629, aes_core_keymem_n628, aes_core_keymem_n627,
         aes_core_keymem_n626, aes_core_keymem_n625, aes_core_keymem_n624,
         aes_core_keymem_n623, aes_core_keymem_n622, aes_core_keymem_n621,
         aes_core_keymem_n620, aes_core_keymem_n619, aes_core_keymem_n618,
         aes_core_keymem_n617, aes_core_keymem_n616, aes_core_keymem_n615,
         aes_core_keymem_n614, aes_core_keymem_n613, aes_core_keymem_n612,
         aes_core_keymem_n611, aes_core_keymem_n610, aes_core_keymem_n609,
         aes_core_keymem_n608, aes_core_keymem_n607, aes_core_keymem_n606,
         aes_core_keymem_n605, aes_core_keymem_n604, aes_core_keymem_n603,
         aes_core_keymem_n602, aes_core_keymem_n601, aes_core_keymem_n600,
         aes_core_keymem_n599, aes_core_keymem_n598, aes_core_keymem_n597,
         aes_core_keymem_n596, aes_core_keymem_n595, aes_core_keymem_n594,
         aes_core_keymem_n593, aes_core_keymem_n592, aes_core_keymem_n591,
         aes_core_keymem_n590, aes_core_keymem_n589, aes_core_keymem_n588,
         aes_core_keymem_n587, aes_core_keymem_n586, aes_core_keymem_n585,
         aes_core_keymem_n584, aes_core_keymem_n583, aes_core_keymem_n582,
         aes_core_keymem_n581, aes_core_keymem_n580, aes_core_keymem_n579,
         aes_core_keymem_n578, aes_core_keymem_n577, aes_core_keymem_n576,
         aes_core_keymem_n575, aes_core_keymem_n574, aes_core_keymem_n573,
         aes_core_keymem_n572, aes_core_keymem_n571, aes_core_keymem_n570,
         aes_core_keymem_n569, aes_core_keymem_n568, aes_core_keymem_n567,
         aes_core_keymem_n566, aes_core_keymem_n565, aes_core_keymem_n564,
         aes_core_keymem_n563, aes_core_keymem_n562, aes_core_keymem_n561,
         aes_core_keymem_n560, aes_core_keymem_n558, aes_core_keymem_n556,
         aes_core_keymem_n555, aes_core_keymem_n553, aes_core_keymem_n552,
         aes_core_keymem_n551, aes_core_keymem_n550, aes_core_keymem_n549,
         aes_core_keymem_n548, aes_core_keymem_n547, aes_core_keymem_n546,
         aes_core_keymem_n545, aes_core_keymem_n543, aes_core_keymem_n542,
         aes_core_keymem_n541, aes_core_keymem_n540, aes_core_keymem_n539,
         aes_core_keymem_n538, aes_core_keymem_n537, aes_core_keymem_n536,
         aes_core_keymem_n535, aes_core_keymem_n534, aes_core_keymem_n533,
         aes_core_keymem_n532, aes_core_keymem_n531, aes_core_keymem_n530,
         aes_core_keymem_n529, aes_core_keymem_n528, aes_core_keymem_n527,
         aes_core_keymem_n526, aes_core_keymem_n525, aes_core_keymem_n524,
         aes_core_keymem_n523, aes_core_keymem_n522, aes_core_keymem_n521,
         aes_core_keymem_n520, aes_core_keymem_n519, aes_core_keymem_n518,
         aes_core_keymem_n517, aes_core_keymem_n516, aes_core_keymem_n515,
         aes_core_keymem_n514, aes_core_keymem_n513, aes_core_keymem_n512,
         aes_core_keymem_n511, aes_core_keymem_n510, aes_core_keymem_n509,
         aes_core_keymem_n508, aes_core_keymem_n507, aes_core_keymem_n506,
         aes_core_keymem_n505, aes_core_keymem_n504, aes_core_keymem_n503,
         aes_core_keymem_n502, aes_core_keymem_n501, aes_core_keymem_n500,
         aes_core_keymem_n499, aes_core_keymem_n498, aes_core_keymem_n497,
         aes_core_keymem_n496, aes_core_keymem_n495, aes_core_keymem_n494,
         aes_core_keymem_n493, aes_core_keymem_n492, aes_core_keymem_n491,
         aes_core_keymem_n490, aes_core_keymem_n489, aes_core_keymem_n488,
         aes_core_keymem_n487, aes_core_keymem_n486, aes_core_keymem_n485,
         aes_core_keymem_n484, aes_core_keymem_n483, aes_core_keymem_n482,
         aes_core_keymem_n481, aes_core_keymem_n480, aes_core_keymem_n479,
         aes_core_keymem_n478, aes_core_keymem_n477, aes_core_keymem_n476,
         aes_core_keymem_n475, aes_core_keymem_n474, aes_core_keymem_n473,
         aes_core_keymem_n472, aes_core_keymem_n471, aes_core_keymem_n470,
         aes_core_keymem_n469, aes_core_keymem_n468, aes_core_keymem_n467,
         aes_core_keymem_n466, aes_core_keymem_n465, aes_core_keymem_n464,
         aes_core_keymem_n463, aes_core_keymem_n462, aes_core_keymem_n461,
         aes_core_keymem_n460, aes_core_keymem_n459, aes_core_keymem_n458,
         aes_core_keymem_n457, aes_core_keymem_n456, aes_core_keymem_n455,
         aes_core_keymem_n454, aes_core_keymem_n453, aes_core_keymem_n452,
         aes_core_keymem_n451, aes_core_keymem_n450, aes_core_keymem_n449,
         aes_core_keymem_n448, aes_core_keymem_n447, aes_core_keymem_n446,
         aes_core_keymem_n445, aes_core_keymem_n444, aes_core_keymem_n443,
         aes_core_keymem_n442, aes_core_keymem_n441, aes_core_keymem_n440,
         aes_core_keymem_n439, aes_core_keymem_n438, aes_core_keymem_n437,
         aes_core_keymem_n436, aes_core_keymem_n435, aes_core_keymem_n434,
         aes_core_keymem_n433, aes_core_keymem_n432, aes_core_keymem_n431,
         aes_core_keymem_n430, aes_core_keymem_n429, aes_core_keymem_n428,
         aes_core_keymem_n427, aes_core_keymem_n426, aes_core_keymem_n425,
         aes_core_keymem_n424, aes_core_keymem_n423, aes_core_keymem_n422,
         aes_core_keymem_n421, aes_core_keymem_n420, aes_core_keymem_n419,
         aes_core_keymem_n418, aes_core_keymem_n417, aes_core_keymem_n416,
         aes_core_keymem_n415, aes_core_keymem_n414, aes_core_keymem_n413,
         aes_core_keymem_n412, aes_core_keymem_n411, aes_core_keymem_n410,
         aes_core_keymem_n409, aes_core_keymem_n408, aes_core_keymem_n407,
         aes_core_keymem_n406, aes_core_keymem_n405, aes_core_keymem_n404,
         aes_core_keymem_n403, aes_core_keymem_n402, aes_core_keymem_n401,
         aes_core_keymem_n400, aes_core_keymem_n399, aes_core_keymem_n398,
         aes_core_keymem_n397, aes_core_keymem_n396, aes_core_keymem_n395,
         aes_core_keymem_n394, aes_core_keymem_n393, aes_core_keymem_n392,
         aes_core_keymem_n391, aes_core_keymem_n390, aes_core_keymem_n389,
         aes_core_keymem_n388, aes_core_keymem_n387, aes_core_keymem_n386,
         aes_core_keymem_n385, aes_core_keymem_n384, aes_core_keymem_n383,
         aes_core_keymem_n382, aes_core_keymem_n381, aes_core_keymem_n380,
         aes_core_keymem_n379, aes_core_keymem_n378, aes_core_keymem_n377,
         aes_core_keymem_n376, aes_core_keymem_n375, aes_core_keymem_n374,
         aes_core_keymem_n373, aes_core_keymem_n372, aes_core_keymem_n371,
         aes_core_keymem_n370, aes_core_keymem_n369, aes_core_keymem_n368,
         aes_core_keymem_n367, aes_core_keymem_n366, aes_core_keymem_n365,
         aes_core_keymem_n364, aes_core_keymem_n363, aes_core_keymem_n362,
         aes_core_keymem_n361, aes_core_keymem_n360, aes_core_keymem_n359,
         aes_core_keymem_n358, aes_core_keymem_n357, aes_core_keymem_n356,
         aes_core_keymem_n355, aes_core_keymem_n354, aes_core_keymem_n353,
         aes_core_keymem_n352, aes_core_keymem_n351, aes_core_keymem_n350,
         aes_core_keymem_n349, aes_core_keymem_n348, aes_core_keymem_n347,
         aes_core_keymem_n346, aes_core_keymem_n345, aes_core_keymem_n344,
         aes_core_keymem_n343, aes_core_keymem_n342, aes_core_keymem_n341,
         aes_core_keymem_n340, aes_core_keymem_n339, aes_core_keymem_n338,
         aes_core_keymem_n337, aes_core_keymem_n336, aes_core_keymem_n335,
         aes_core_keymem_n334, aes_core_keymem_n333, aes_core_keymem_n332,
         aes_core_keymem_n331, aes_core_keymem_n330, aes_core_keymem_n329,
         aes_core_keymem_n328, aes_core_keymem_n327, aes_core_keymem_n326,
         aes_core_keymem_n325, aes_core_keymem_n324, aes_core_keymem_n323,
         aes_core_keymem_n322, aes_core_keymem_n321, aes_core_keymem_n320,
         aes_core_keymem_n319, aes_core_keymem_n318, aes_core_keymem_n317,
         aes_core_keymem_n316, aes_core_keymem_n315, aes_core_keymem_n314,
         aes_core_keymem_n313, aes_core_keymem_n312, aes_core_keymem_n311,
         aes_core_keymem_n310, aes_core_keymem_n309, aes_core_keymem_n308,
         aes_core_keymem_n307, aes_core_keymem_n306, aes_core_keymem_n305,
         aes_core_keymem_n304, aes_core_keymem_n303, aes_core_keymem_n302,
         aes_core_keymem_n301, aes_core_keymem_n300, aes_core_keymem_n299,
         aes_core_keymem_n298, aes_core_keymem_n297, aes_core_keymem_n296,
         aes_core_keymem_n295, aes_core_keymem_n294, aes_core_keymem_n293,
         aes_core_keymem_n292, aes_core_keymem_n291, aes_core_keymem_n290,
         aes_core_keymem_n289, aes_core_keymem_n288, aes_core_keymem_n287,
         aes_core_keymem_n286, aes_core_keymem_n285, aes_core_keymem_n284,
         aes_core_keymem_n283, aes_core_keymem_n282, aes_core_keymem_n281,
         aes_core_keymem_n280, aes_core_keymem_n279, aes_core_keymem_n278,
         aes_core_keymem_n277, aes_core_keymem_n276, aes_core_keymem_n275,
         aes_core_keymem_n274, aes_core_keymem_n273, aes_core_keymem_n272,
         aes_core_keymem_n271, aes_core_keymem_n270, aes_core_keymem_n269,
         aes_core_keymem_n268, aes_core_keymem_n267, aes_core_keymem_n266,
         aes_core_keymem_n265, aes_core_keymem_n264, aes_core_keymem_n263,
         aes_core_keymem_n262, aes_core_keymem_n261, aes_core_keymem_n260,
         aes_core_keymem_n259, aes_core_keymem_n258, aes_core_keymem_n257,
         aes_core_keymem_n256, aes_core_keymem_n255, aes_core_keymem_n254,
         aes_core_keymem_n253, aes_core_keymem_n252, aes_core_keymem_n251,
         aes_core_keymem_n250, aes_core_keymem_n249, aes_core_keymem_n248,
         aes_core_keymem_n247, aes_core_keymem_n246, aes_core_keymem_n245,
         aes_core_keymem_n244, aes_core_keymem_n243, aes_core_keymem_n242,
         aes_core_keymem_n241, aes_core_keymem_n240, aes_core_keymem_n239,
         aes_core_keymem_n238, aes_core_keymem_n237, aes_core_keymem_n236,
         aes_core_keymem_n235, aes_core_keymem_n234, aes_core_keymem_n233,
         aes_core_keymem_n232, aes_core_keymem_n231, aes_core_keymem_n230,
         aes_core_keymem_n229, aes_core_keymem_n228, aes_core_keymem_n227,
         aes_core_keymem_n226, aes_core_keymem_n225, aes_core_keymem_n224,
         aes_core_keymem_n223, aes_core_keymem_n222, aes_core_keymem_n221,
         aes_core_keymem_n220, aes_core_keymem_n219, aes_core_keymem_n218,
         aes_core_keymem_n217, aes_core_keymem_n216, aes_core_keymem_n215,
         aes_core_keymem_n214, aes_core_keymem_n213, aes_core_keymem_n212,
         aes_core_keymem_n211, aes_core_keymem_n210, aes_core_keymem_n209,
         aes_core_keymem_n208, aes_core_keymem_n207, aes_core_keymem_n206,
         aes_core_keymem_n205, aes_core_keymem_n204, aes_core_keymem_n203,
         aes_core_keymem_n202, aes_core_keymem_n201, aes_core_keymem_n200,
         aes_core_keymem_n199, aes_core_keymem_n198, aes_core_keymem_n197,
         aes_core_keymem_n196, aes_core_keymem_n195, aes_core_keymem_n194,
         aes_core_keymem_n193, aes_core_keymem_n192, aes_core_keymem_n191,
         aes_core_keymem_n190, aes_core_keymem_n189, aes_core_keymem_n188,
         aes_core_keymem_n187, aes_core_keymem_n186, aes_core_keymem_n185,
         aes_core_keymem_n184, aes_core_keymem_n183, aes_core_keymem_n182,
         aes_core_keymem_n181, aes_core_keymem_n180, aes_core_keymem_n179,
         aes_core_keymem_n178, aes_core_keymem_n177, aes_core_keymem_n176,
         aes_core_keymem_n175, aes_core_keymem_n174, aes_core_keymem_n173,
         aes_core_keymem_n172, aes_core_keymem_n171, aes_core_keymem_n170,
         aes_core_keymem_n169, aes_core_keymem_n168, aes_core_keymem_n167,
         aes_core_keymem_n166, aes_core_keymem_n165, aes_core_keymem_n164,
         aes_core_keymem_n163, aes_core_keymem_n162, aes_core_keymem_n161,
         aes_core_keymem_n160, aes_core_keymem_n159, aes_core_keymem_n158,
         aes_core_keymem_n157, aes_core_keymem_n156, aes_core_keymem_n155,
         aes_core_keymem_n154, aes_core_keymem_n153, aes_core_keymem_n152,
         aes_core_keymem_n151, aes_core_keymem_n150, aes_core_keymem_n149,
         aes_core_keymem_n148, aes_core_keymem_n147, aes_core_keymem_n146,
         aes_core_keymem_n145, aes_core_keymem_n144, aes_core_keymem_n143,
         aes_core_keymem_n142, aes_core_keymem_n141, aes_core_keymem_n140,
         aes_core_keymem_n139, aes_core_keymem_n138, aes_core_keymem_n137,
         aes_core_keymem_n136, aes_core_keymem_n135, aes_core_keymem_n134,
         aes_core_keymem_n133, aes_core_keymem_n132, aes_core_keymem_n131,
         aes_core_keymem_n130, aes_core_keymem_n129, aes_core_keymem_n128,
         aes_core_keymem_n127, aes_core_keymem_n126, aes_core_keymem_n125,
         aes_core_keymem_n124, aes_core_keymem_n123, aes_core_keymem_n122,
         aes_core_keymem_n121, aes_core_keymem_n120, aes_core_keymem_n119,
         aes_core_keymem_n118, aes_core_keymem_n117, aes_core_keymem_n116,
         aes_core_keymem_n115, aes_core_keymem_n114, aes_core_keymem_n113,
         aes_core_keymem_n112, aes_core_keymem_n111, aes_core_keymem_n110,
         aes_core_keymem_n109, aes_core_keymem_n108, aes_core_keymem_n107,
         aes_core_keymem_n106, aes_core_keymem_n105, aes_core_keymem_n104,
         aes_core_keymem_n103, aes_core_keymem_n102, aes_core_keymem_n101,
         aes_core_keymem_n100, aes_core_keymem_n99, aes_core_keymem_n98,
         aes_core_keymem_n97, aes_core_keymem_n96, aes_core_keymem_n95,
         aes_core_keymem_n94, aes_core_keymem_n93, aes_core_keymem_n92,
         aes_core_keymem_n91, aes_core_keymem_n90, aes_core_keymem_n89,
         aes_core_keymem_n88, aes_core_keymem_n87, aes_core_keymem_n86,
         aes_core_keymem_n85, aes_core_keymem_n84, aes_core_keymem_n83,
         aes_core_keymem_n82, aes_core_keymem_n81, aes_core_keymem_n80,
         aes_core_keymem_n79, aes_core_keymem_n78, aes_core_keymem_n77,
         aes_core_keymem_n76, aes_core_keymem_n75, aes_core_keymem_n74,
         aes_core_keymem_n73, aes_core_keymem_n72, aes_core_keymem_n71,
         aes_core_keymem_n70, aes_core_keymem_n69, aes_core_keymem_n68,
         aes_core_keymem_n67, aes_core_keymem_n66, aes_core_keymem_n65,
         aes_core_keymem_n64, aes_core_keymem_n63, aes_core_keymem_n62,
         aes_core_keymem_n61, aes_core_keymem_n60, aes_core_keymem_n59,
         aes_core_keymem_n58, aes_core_keymem_n57, aes_core_keymem_n56,
         aes_core_keymem_n55, aes_core_keymem_n54, aes_core_keymem_n53,
         aes_core_keymem_n52, aes_core_keymem_n51, aes_core_keymem_n50,
         aes_core_keymem_n49, aes_core_keymem_n48, aes_core_keymem_n47,
         aes_core_keymem_n46, aes_core_keymem_n45, aes_core_keymem_n44,
         aes_core_keymem_n43, aes_core_keymem_n42, aes_core_keymem_n41,
         aes_core_keymem_n40, aes_core_keymem_n39, aes_core_keymem_n38,
         aes_core_keymem_n37, aes_core_keymem_n36, aes_core_keymem_n35,
         aes_core_keymem_n34, aes_core_keymem_n33, aes_core_keymem_n32,
         aes_core_keymem_n31, aes_core_keymem_n29, aes_core_keymem_n28,
         aes_core_keymem_n27, aes_core_keymem_n26, aes_core_keymem_n25,
         aes_core_keymem_n23, aes_core_keymem_n21, aes_core_keymem_n20,
         aes_core_keymem_n19, aes_core_keymem_n18, aes_core_keymem_n14,
         aes_core_keymem_n9, aes_core_sbox_inst_n1735,
         aes_core_sbox_inst_n1734, aes_core_sbox_inst_n1733,
         aes_core_sbox_inst_n1732, aes_core_sbox_inst_n1731,
         aes_core_sbox_inst_n1730, aes_core_sbox_inst_n1729,
         aes_core_sbox_inst_n1728, aes_core_sbox_inst_n1727,
         aes_core_sbox_inst_n1726, aes_core_sbox_inst_n1725,
         aes_core_sbox_inst_n1724, aes_core_sbox_inst_n1723,
         aes_core_sbox_inst_n1722, aes_core_sbox_inst_n1721,
         aes_core_sbox_inst_n1720, aes_core_sbox_inst_n1719,
         aes_core_sbox_inst_n1718, aes_core_sbox_inst_n1717,
         aes_core_sbox_inst_n1716, aes_core_sbox_inst_n1715,
         aes_core_sbox_inst_n1714, aes_core_sbox_inst_n1713,
         aes_core_sbox_inst_n1712, aes_core_sbox_inst_n1711,
         aes_core_sbox_inst_n1710, aes_core_sbox_inst_n1709,
         aes_core_sbox_inst_n1708, aes_core_sbox_inst_n1707,
         aes_core_sbox_inst_n1706, aes_core_sbox_inst_n1705,
         aes_core_sbox_inst_n1704, aes_core_sbox_inst_n1703,
         aes_core_sbox_inst_n1702, aes_core_sbox_inst_n1701,
         aes_core_sbox_inst_n1700, aes_core_sbox_inst_n1699,
         aes_core_sbox_inst_n1698, aes_core_sbox_inst_n1697,
         aes_core_sbox_inst_n1696, aes_core_sbox_inst_n1695,
         aes_core_sbox_inst_n1694, aes_core_sbox_inst_n1693,
         aes_core_sbox_inst_n1692, aes_core_sbox_inst_n1691,
         aes_core_sbox_inst_n1690, aes_core_sbox_inst_n1689,
         aes_core_sbox_inst_n1688, aes_core_sbox_inst_n1687,
         aes_core_sbox_inst_n1686, aes_core_sbox_inst_n1685,
         aes_core_sbox_inst_n1684, aes_core_sbox_inst_n1683,
         aes_core_sbox_inst_n1682, aes_core_sbox_inst_n1681,
         aes_core_sbox_inst_n1680, aes_core_sbox_inst_n1679,
         aes_core_sbox_inst_n1678, aes_core_sbox_inst_n1677,
         aes_core_sbox_inst_n1676, aes_core_sbox_inst_n1675,
         aes_core_sbox_inst_n1674, aes_core_sbox_inst_n1673,
         aes_core_sbox_inst_n1672, aes_core_sbox_inst_n1671,
         aes_core_sbox_inst_n1670, aes_core_sbox_inst_n1669,
         aes_core_sbox_inst_n1668, aes_core_sbox_inst_n1667,
         aes_core_sbox_inst_n1666, aes_core_sbox_inst_n1665,
         aes_core_sbox_inst_n1664, aes_core_sbox_inst_n1663,
         aes_core_sbox_inst_n1662, aes_core_sbox_inst_n1661,
         aes_core_sbox_inst_n1660, aes_core_sbox_inst_n1659,
         aes_core_sbox_inst_n1658, aes_core_sbox_inst_n1657,
         aes_core_sbox_inst_n1656, aes_core_sbox_inst_n1655,
         aes_core_sbox_inst_n1654, aes_core_sbox_inst_n1653,
         aes_core_sbox_inst_n1652, aes_core_sbox_inst_n1651,
         aes_core_sbox_inst_n1650, aes_core_sbox_inst_n1649,
         aes_core_sbox_inst_n1648, aes_core_sbox_inst_n1647,
         aes_core_sbox_inst_n1646, aes_core_sbox_inst_n1645,
         aes_core_sbox_inst_n1644, aes_core_sbox_inst_n1643,
         aes_core_sbox_inst_n1642, aes_core_sbox_inst_n1641,
         aes_core_sbox_inst_n1640, aes_core_sbox_inst_n1639,
         aes_core_sbox_inst_n1638, aes_core_sbox_inst_n1637,
         aes_core_sbox_inst_n1636, aes_core_sbox_inst_n1635,
         aes_core_sbox_inst_n1634, aes_core_sbox_inst_n1633,
         aes_core_sbox_inst_n1632, aes_core_sbox_inst_n1631,
         aes_core_sbox_inst_n1630, aes_core_sbox_inst_n1629,
         aes_core_sbox_inst_n1628, aes_core_sbox_inst_n1627,
         aes_core_sbox_inst_n1626, aes_core_sbox_inst_n1625,
         aes_core_sbox_inst_n1624, aes_core_sbox_inst_n1623,
         aes_core_sbox_inst_n1622, aes_core_sbox_inst_n1621,
         aes_core_sbox_inst_n1620, aes_core_sbox_inst_n1619,
         aes_core_sbox_inst_n1618, aes_core_sbox_inst_n1617,
         aes_core_sbox_inst_n1616, aes_core_sbox_inst_n1615,
         aes_core_sbox_inst_n1614, aes_core_sbox_inst_n1613,
         aes_core_sbox_inst_n1612, aes_core_sbox_inst_n1611,
         aes_core_sbox_inst_n1610, aes_core_sbox_inst_n1609,
         aes_core_sbox_inst_n1608, aes_core_sbox_inst_n1607,
         aes_core_sbox_inst_n1606, aes_core_sbox_inst_n1605,
         aes_core_sbox_inst_n1604, aes_core_sbox_inst_n1603,
         aes_core_sbox_inst_n1602, aes_core_sbox_inst_n1601,
         aes_core_sbox_inst_n1600, aes_core_sbox_inst_n1599,
         aes_core_sbox_inst_n1598, aes_core_sbox_inst_n1597,
         aes_core_sbox_inst_n1596, aes_core_sbox_inst_n1595,
         aes_core_sbox_inst_n1594, aes_core_sbox_inst_n1593,
         aes_core_sbox_inst_n1592, aes_core_sbox_inst_n1591,
         aes_core_sbox_inst_n1590, aes_core_sbox_inst_n1589,
         aes_core_sbox_inst_n1588, aes_core_sbox_inst_n1587,
         aes_core_sbox_inst_n1586, aes_core_sbox_inst_n1585,
         aes_core_sbox_inst_n1584, aes_core_sbox_inst_n1583,
         aes_core_sbox_inst_n1582, aes_core_sbox_inst_n1581,
         aes_core_sbox_inst_n1580, aes_core_sbox_inst_n1579,
         aes_core_sbox_inst_n1578, aes_core_sbox_inst_n1577,
         aes_core_sbox_inst_n1576, aes_core_sbox_inst_n1575,
         aes_core_sbox_inst_n1574, aes_core_sbox_inst_n1573,
         aes_core_sbox_inst_n1572, aes_core_sbox_inst_n1571,
         aes_core_sbox_inst_n1570, aes_core_sbox_inst_n1569,
         aes_core_sbox_inst_n1568, aes_core_sbox_inst_n1567,
         aes_core_sbox_inst_n1566, aes_core_sbox_inst_n617,
         aes_core_sbox_inst_n450, aes_core_sbox_inst_n316,
         aes_core_sbox_inst_n273, aes_core_sbox_inst_n259,
         aes_core_sbox_inst_n258, aes_core_sbox_inst_n257,
         aes_core_sbox_inst_n256, aes_core_sbox_inst_n255,
         aes_core_sbox_inst_n254, aes_core_sbox_inst_n253,
         aes_core_sbox_inst_n252, aes_core_sbox_inst_n251,
         aes_core_sbox_inst_n250, aes_core_sbox_inst_n249,
         aes_core_sbox_inst_n248, aes_core_sbox_inst_n247,
         aes_core_sbox_inst_n246, aes_core_sbox_inst_n245,
         aes_core_sbox_inst_n244, aes_core_sbox_inst_n243,
         aes_core_sbox_inst_n242, aes_core_sbox_inst_n241,
         aes_core_sbox_inst_n240, aes_core_sbox_inst_n239,
         aes_core_sbox_inst_n238, aes_core_sbox_inst_n237,
         aes_core_sbox_inst_n236, aes_core_sbox_inst_n235,
         aes_core_sbox_inst_n234, aes_core_sbox_inst_n233,
         aes_core_sbox_inst_n232, aes_core_sbox_inst_n231,
         aes_core_sbox_inst_n230, aes_core_sbox_inst_n229,
         aes_core_sbox_inst_n228, aes_core_sbox_inst_n227,
         aes_core_sbox_inst_n226, aes_core_sbox_inst_n225,
         aes_core_sbox_inst_n224, aes_core_sbox_inst_n223,
         aes_core_sbox_inst_n222, aes_core_sbox_inst_n221,
         aes_core_sbox_inst_n220, aes_core_sbox_inst_n219,
         aes_core_sbox_inst_n218, aes_core_sbox_inst_n217,
         aes_core_sbox_inst_n216, aes_core_sbox_inst_n215,
         aes_core_sbox_inst_n214, aes_core_sbox_inst_n213,
         aes_core_sbox_inst_n212, aes_core_sbox_inst_n211,
         aes_core_sbox_inst_n210, aes_core_sbox_inst_n209,
         aes_core_sbox_inst_n208, aes_core_sbox_inst_n207,
         aes_core_sbox_inst_n206, aes_core_sbox_inst_n205,
         aes_core_sbox_inst_n204, aes_core_sbox_inst_n203,
         aes_core_sbox_inst_n202, aes_core_sbox_inst_n201,
         aes_core_sbox_inst_n200, aes_core_sbox_inst_n199,
         aes_core_sbox_inst_n198, aes_core_sbox_inst_n197,
         aes_core_sbox_inst_n196, aes_core_sbox_inst_n195,
         aes_core_sbox_inst_n194, aes_core_sbox_inst_n193,
         aes_core_sbox_inst_n192, aes_core_sbox_inst_n191,
         aes_core_sbox_inst_n190, aes_core_sbox_inst_n189,
         aes_core_sbox_inst_n188, aes_core_sbox_inst_n187,
         aes_core_sbox_inst_n186, aes_core_sbox_inst_n185,
         aes_core_sbox_inst_n184, aes_core_sbox_inst_n183,
         aes_core_sbox_inst_n182, aes_core_sbox_inst_n181,
         aes_core_sbox_inst_n180, aes_core_sbox_inst_n179,
         aes_core_sbox_inst_n178, aes_core_sbox_inst_n177,
         aes_core_sbox_inst_n176, aes_core_sbox_inst_n175,
         aes_core_sbox_inst_n174, aes_core_sbox_inst_n173,
         aes_core_sbox_inst_n172, aes_core_sbox_inst_n171,
         aes_core_sbox_inst_n170, aes_core_sbox_inst_n169,
         aes_core_sbox_inst_n168, aes_core_sbox_inst_n167,
         aes_core_sbox_inst_n166, aes_core_sbox_inst_n165,
         aes_core_sbox_inst_n164, aes_core_sbox_inst_n163,
         aes_core_sbox_inst_n162, aes_core_sbox_inst_n161,
         aes_core_sbox_inst_n160, aes_core_sbox_inst_n159,
         aes_core_sbox_inst_n158, aes_core_sbox_inst_n157,
         aes_core_sbox_inst_n156, aes_core_sbox_inst_n155,
         aes_core_sbox_inst_n154, aes_core_sbox_inst_n153,
         aes_core_sbox_inst_n152, aes_core_sbox_inst_n151,
         aes_core_sbox_inst_n150, aes_core_sbox_inst_n149,
         aes_core_sbox_inst_n148, aes_core_sbox_inst_n147,
         aes_core_sbox_inst_n146, aes_core_sbox_inst_n145,
         aes_core_sbox_inst_n144, aes_core_sbox_inst_n143,
         aes_core_sbox_inst_n142, aes_core_sbox_inst_n141,
         aes_core_sbox_inst_n140, aes_core_sbox_inst_n139,
         aes_core_sbox_inst_n138, aes_core_sbox_inst_n137,
         aes_core_sbox_inst_n136, aes_core_sbox_inst_n135,
         aes_core_sbox_inst_n134, aes_core_sbox_inst_n133,
         aes_core_sbox_inst_n132, aes_core_sbox_inst_n131,
         aes_core_sbox_inst_n130, aes_core_sbox_inst_n129,
         aes_core_sbox_inst_n128, aes_core_sbox_inst_n127,
         aes_core_sbox_inst_n126, aes_core_sbox_inst_n125,
         aes_core_sbox_inst_n124, aes_core_sbox_inst_n123,
         aes_core_sbox_inst_n122, aes_core_sbox_inst_n121,
         aes_core_sbox_inst_n120, aes_core_sbox_inst_n119,
         aes_core_sbox_inst_n118, aes_core_sbox_inst_n117,
         aes_core_sbox_inst_n116, aes_core_sbox_inst_n115,
         aes_core_sbox_inst_n114, aes_core_sbox_inst_n113,
         aes_core_sbox_inst_n112, aes_core_sbox_inst_n111,
         aes_core_sbox_inst_n110, aes_core_sbox_inst_n109,
         aes_core_sbox_inst_n108, aes_core_sbox_inst_n107,
         aes_core_sbox_inst_n106, aes_core_sbox_inst_n105,
         aes_core_sbox_inst_n104, aes_core_sbox_inst_n103,
         aes_core_sbox_inst_n102, aes_core_sbox_inst_n101,
         aes_core_sbox_inst_n100, aes_core_sbox_inst_n99,
         aes_core_sbox_inst_n98, aes_core_sbox_inst_n97,
         aes_core_sbox_inst_n96, aes_core_sbox_inst_n95,
         aes_core_sbox_inst_n94, aes_core_sbox_inst_n93,
         aes_core_sbox_inst_n92, aes_core_sbox_inst_n91,
         aes_core_sbox_inst_n90, aes_core_sbox_inst_n89,
         aes_core_sbox_inst_n88, aes_core_sbox_inst_n87,
         aes_core_sbox_inst_n86, aes_core_sbox_inst_n85,
         aes_core_sbox_inst_n84, aes_core_sbox_inst_n83,
         aes_core_sbox_inst_n82, aes_core_sbox_inst_n81,
         aes_core_sbox_inst_n80, aes_core_sbox_inst_n79,
         aes_core_sbox_inst_n78, aes_core_sbox_inst_n77,
         aes_core_sbox_inst_n76, aes_core_sbox_inst_n75,
         aes_core_sbox_inst_n74, aes_core_sbox_inst_n73,
         aes_core_sbox_inst_n72, aes_core_sbox_inst_n71,
         aes_core_sbox_inst_n70, aes_core_sbox_inst_n69,
         aes_core_sbox_inst_n68, aes_core_sbox_inst_n67,
         aes_core_sbox_inst_n66, aes_core_sbox_inst_n65,
         aes_core_sbox_inst_n64, aes_core_sbox_inst_n63,
         aes_core_sbox_inst_n62, aes_core_sbox_inst_n61,
         aes_core_sbox_inst_n60, aes_core_sbox_inst_n59,
         aes_core_sbox_inst_n58, aes_core_sbox_inst_n57,
         aes_core_sbox_inst_n56, aes_core_sbox_inst_n55,
         aes_core_sbox_inst_n54, aes_core_sbox_inst_n53,
         aes_core_sbox_inst_n52, aes_core_sbox_inst_n51,
         aes_core_sbox_inst_n50, aes_core_sbox_inst_n49,
         aes_core_sbox_inst_n48, aes_core_sbox_inst_n47,
         aes_core_sbox_inst_n46, aes_core_sbox_inst_n45,
         aes_core_sbox_inst_n44, aes_core_sbox_inst_n43,
         aes_core_sbox_inst_n42, aes_core_sbox_inst_n41,
         aes_core_sbox_inst_n40, aes_core_sbox_inst_n39,
         aes_core_sbox_inst_n38, aes_core_sbox_inst_n37,
         aes_core_sbox_inst_n36, aes_core_sbox_inst_n35,
         aes_core_sbox_inst_n34, aes_core_sbox_inst_n33,
         aes_core_sbox_inst_n32, aes_core_sbox_inst_n31,
         aes_core_sbox_inst_n30, aes_core_sbox_inst_n29,
         aes_core_sbox_inst_n28, aes_core_sbox_inst_n27,
         aes_core_sbox_inst_n26, aes_core_sbox_inst_n25,
         aes_core_sbox_inst_n24, aes_core_sbox_inst_n23,
         aes_core_sbox_inst_n22, aes_core_sbox_inst_n21,
         aes_core_sbox_inst_n20, aes_core_sbox_inst_n19,
         aes_core_sbox_inst_n18, aes_core_sbox_inst_n17,
         aes_core_sbox_inst_n16, aes_core_sbox_inst_n15,
         aes_core_sbox_inst_n14, aes_core_sbox_inst_n13,
         aes_core_sbox_inst_n12, aes_core_sbox_inst_n11,
         aes_core_sbox_inst_n10, aes_core_sbox_inst_n9, aes_core_sbox_inst_n8,
         aes_core_sbox_inst_n7, aes_core_sbox_inst_n6, aes_core_sbox_inst_n5,
         aes_core_sbox_inst_n4, aes_core_sbox_inst_n3, aes_core_sbox_inst_n2,
         aes_core_sbox_inst_n1, aes_core_sbox_inst_n1565,
         aes_core_sbox_inst_n1564, aes_core_sbox_inst_n1563,
         aes_core_sbox_inst_n1562, aes_core_sbox_inst_n1561,
         aes_core_sbox_inst_n1560, aes_core_sbox_inst_n1559,
         aes_core_sbox_inst_n1558, aes_core_sbox_inst_n1557,
         aes_core_sbox_inst_n1556, aes_core_sbox_inst_n1555,
         aes_core_sbox_inst_n1554, aes_core_sbox_inst_n1553,
         aes_core_sbox_inst_n1552, aes_core_sbox_inst_n1551,
         aes_core_sbox_inst_n1550, aes_core_sbox_inst_n1549,
         aes_core_sbox_inst_n1548, aes_core_sbox_inst_n1547,
         aes_core_sbox_inst_n1546, aes_core_sbox_inst_n1545,
         aes_core_sbox_inst_n1544, aes_core_sbox_inst_n1543,
         aes_core_sbox_inst_n1542, aes_core_sbox_inst_n1541,
         aes_core_sbox_inst_n1540, aes_core_sbox_inst_n1539,
         aes_core_sbox_inst_n1538, aes_core_sbox_inst_n1537,
         aes_core_sbox_inst_n1536, aes_core_sbox_inst_n1535,
         aes_core_sbox_inst_n1534, aes_core_sbox_inst_n1533,
         aes_core_sbox_inst_n1532, aes_core_sbox_inst_n1531,
         aes_core_sbox_inst_n1530, aes_core_sbox_inst_n1529,
         aes_core_sbox_inst_n1528, aes_core_sbox_inst_n1527,
         aes_core_sbox_inst_n1526, aes_core_sbox_inst_n1525,
         aes_core_sbox_inst_n1524, aes_core_sbox_inst_n1523,
         aes_core_sbox_inst_n1522, aes_core_sbox_inst_n1521,
         aes_core_sbox_inst_n1520, aes_core_sbox_inst_n1519,
         aes_core_sbox_inst_n1518, aes_core_sbox_inst_n1517,
         aes_core_sbox_inst_n1516, aes_core_sbox_inst_n1515,
         aes_core_sbox_inst_n1514, aes_core_sbox_inst_n1513,
         aes_core_sbox_inst_n1512, aes_core_sbox_inst_n1511,
         aes_core_sbox_inst_n1510, aes_core_sbox_inst_n1509,
         aes_core_sbox_inst_n1508, aes_core_sbox_inst_n1507,
         aes_core_sbox_inst_n1506, aes_core_sbox_inst_n1505,
         aes_core_sbox_inst_n1504, aes_core_sbox_inst_n1503,
         aes_core_sbox_inst_n1502, aes_core_sbox_inst_n1501,
         aes_core_sbox_inst_n1500, aes_core_sbox_inst_n1499,
         aes_core_sbox_inst_n1498, aes_core_sbox_inst_n1497,
         aes_core_sbox_inst_n1496, aes_core_sbox_inst_n1495,
         aes_core_sbox_inst_n1494, aes_core_sbox_inst_n1493,
         aes_core_sbox_inst_n1492, aes_core_sbox_inst_n1491,
         aes_core_sbox_inst_n1490, aes_core_sbox_inst_n1489,
         aes_core_sbox_inst_n1488, aes_core_sbox_inst_n1487,
         aes_core_sbox_inst_n1486, aes_core_sbox_inst_n1485,
         aes_core_sbox_inst_n1484, aes_core_sbox_inst_n1483,
         aes_core_sbox_inst_n1482, aes_core_sbox_inst_n1481,
         aes_core_sbox_inst_n1480, aes_core_sbox_inst_n1479,
         aes_core_sbox_inst_n1478, aes_core_sbox_inst_n1477,
         aes_core_sbox_inst_n1476, aes_core_sbox_inst_n1475,
         aes_core_sbox_inst_n1474, aes_core_sbox_inst_n1473,
         aes_core_sbox_inst_n1472, aes_core_sbox_inst_n1471,
         aes_core_sbox_inst_n1470, aes_core_sbox_inst_n1469,
         aes_core_sbox_inst_n1468, aes_core_sbox_inst_n1467,
         aes_core_sbox_inst_n1466, aes_core_sbox_inst_n1465,
         aes_core_sbox_inst_n1464, aes_core_sbox_inst_n1463,
         aes_core_sbox_inst_n1462, aes_core_sbox_inst_n1461,
         aes_core_sbox_inst_n1460, aes_core_sbox_inst_n1459,
         aes_core_sbox_inst_n1458, aes_core_sbox_inst_n1457,
         aes_core_sbox_inst_n1456, aes_core_sbox_inst_n1455,
         aes_core_sbox_inst_n1454, aes_core_sbox_inst_n1453,
         aes_core_sbox_inst_n1452, aes_core_sbox_inst_n1451,
         aes_core_sbox_inst_n1450, aes_core_sbox_inst_n1449,
         aes_core_sbox_inst_n1448, aes_core_sbox_inst_n1447,
         aes_core_sbox_inst_n1446, aes_core_sbox_inst_n1445,
         aes_core_sbox_inst_n1444, aes_core_sbox_inst_n1443,
         aes_core_sbox_inst_n1442, aes_core_sbox_inst_n1441,
         aes_core_sbox_inst_n1440, aes_core_sbox_inst_n1439,
         aes_core_sbox_inst_n1438, aes_core_sbox_inst_n1437,
         aes_core_sbox_inst_n1436, aes_core_sbox_inst_n1435,
         aes_core_sbox_inst_n1434, aes_core_sbox_inst_n1433,
         aes_core_sbox_inst_n1432, aes_core_sbox_inst_n1431,
         aes_core_sbox_inst_n1430, aes_core_sbox_inst_n1429,
         aes_core_sbox_inst_n1428, aes_core_sbox_inst_n1427,
         aes_core_sbox_inst_n1426, aes_core_sbox_inst_n1425,
         aes_core_sbox_inst_n1424, aes_core_sbox_inst_n1423,
         aes_core_sbox_inst_n1422, aes_core_sbox_inst_n1421,
         aes_core_sbox_inst_n1420, aes_core_sbox_inst_n1419,
         aes_core_sbox_inst_n1418, aes_core_sbox_inst_n1417,
         aes_core_sbox_inst_n1416, aes_core_sbox_inst_n1415,
         aes_core_sbox_inst_n1414, aes_core_sbox_inst_n1413,
         aes_core_sbox_inst_n1412, aes_core_sbox_inst_n1411,
         aes_core_sbox_inst_n1410, aes_core_sbox_inst_n1409,
         aes_core_sbox_inst_n1408, aes_core_sbox_inst_n1407,
         aes_core_sbox_inst_n1406, aes_core_sbox_inst_n1405,
         aes_core_sbox_inst_n1404, aes_core_sbox_inst_n1403,
         aes_core_sbox_inst_n1402, aes_core_sbox_inst_n1401,
         aes_core_sbox_inst_n1400, aes_core_sbox_inst_n1399,
         aes_core_sbox_inst_n1398, aes_core_sbox_inst_n1397,
         aes_core_sbox_inst_n1396, aes_core_sbox_inst_n1395,
         aes_core_sbox_inst_n1394, aes_core_sbox_inst_n1393,
         aes_core_sbox_inst_n1392, aes_core_sbox_inst_n1391,
         aes_core_sbox_inst_n1390, aes_core_sbox_inst_n1389,
         aes_core_sbox_inst_n1388, aes_core_sbox_inst_n1387,
         aes_core_sbox_inst_n1386, aes_core_sbox_inst_n1385,
         aes_core_sbox_inst_n1384, aes_core_sbox_inst_n1383,
         aes_core_sbox_inst_n1382, aes_core_sbox_inst_n1381,
         aes_core_sbox_inst_n1380, aes_core_sbox_inst_n1379,
         aes_core_sbox_inst_n1378, aes_core_sbox_inst_n1377,
         aes_core_sbox_inst_n1376, aes_core_sbox_inst_n1375,
         aes_core_sbox_inst_n1374, aes_core_sbox_inst_n1373,
         aes_core_sbox_inst_n1372, aes_core_sbox_inst_n1371,
         aes_core_sbox_inst_n1370, aes_core_sbox_inst_n1369,
         aes_core_sbox_inst_n1368, aes_core_sbox_inst_n1367,
         aes_core_sbox_inst_n1366, aes_core_sbox_inst_n1365,
         aes_core_sbox_inst_n1364, aes_core_sbox_inst_n1363,
         aes_core_sbox_inst_n1362, aes_core_sbox_inst_n1361,
         aes_core_sbox_inst_n1360, aes_core_sbox_inst_n1359,
         aes_core_sbox_inst_n1358, aes_core_sbox_inst_n1357,
         aes_core_sbox_inst_n1356, aes_core_sbox_inst_n1355,
         aes_core_sbox_inst_n1354, aes_core_sbox_inst_n1353,
         aes_core_sbox_inst_n1352, aes_core_sbox_inst_n1351,
         aes_core_sbox_inst_n1350, aes_core_sbox_inst_n1349,
         aes_core_sbox_inst_n1348, aes_core_sbox_inst_n1347,
         aes_core_sbox_inst_n1346, aes_core_sbox_inst_n1345,
         aes_core_sbox_inst_n1344, aes_core_sbox_inst_n1343,
         aes_core_sbox_inst_n1342, aes_core_sbox_inst_n1341,
         aes_core_sbox_inst_n1340, aes_core_sbox_inst_n1339,
         aes_core_sbox_inst_n1338, aes_core_sbox_inst_n1337,
         aes_core_sbox_inst_n1336, aes_core_sbox_inst_n1335,
         aes_core_sbox_inst_n1334, aes_core_sbox_inst_n1333,
         aes_core_sbox_inst_n1332, aes_core_sbox_inst_n1331,
         aes_core_sbox_inst_n1330, aes_core_sbox_inst_n1329,
         aes_core_sbox_inst_n1328, aes_core_sbox_inst_n1327,
         aes_core_sbox_inst_n1326, aes_core_sbox_inst_n1325,
         aes_core_sbox_inst_n1324, aes_core_sbox_inst_n1323,
         aes_core_sbox_inst_n1322, aes_core_sbox_inst_n1321,
         aes_core_sbox_inst_n1320, aes_core_sbox_inst_n1319,
         aes_core_sbox_inst_n1318, aes_core_sbox_inst_n1317,
         aes_core_sbox_inst_n1316, aes_core_sbox_inst_n1315,
         aes_core_sbox_inst_n1314, aes_core_sbox_inst_n1313,
         aes_core_sbox_inst_n1312, aes_core_sbox_inst_n1311,
         aes_core_sbox_inst_n1310, aes_core_sbox_inst_n1309,
         aes_core_sbox_inst_n1308, aes_core_sbox_inst_n1307,
         aes_core_sbox_inst_n1306, aes_core_sbox_inst_n1305,
         aes_core_sbox_inst_n1304, aes_core_sbox_inst_n1303,
         aes_core_sbox_inst_n1302, aes_core_sbox_inst_n1301,
         aes_core_sbox_inst_n1300, aes_core_sbox_inst_n1299,
         aes_core_sbox_inst_n1298, aes_core_sbox_inst_n1297,
         aes_core_sbox_inst_n1296, aes_core_sbox_inst_n1295,
         aes_core_sbox_inst_n1294, aes_core_sbox_inst_n1293,
         aes_core_sbox_inst_n1292, aes_core_sbox_inst_n1291,
         aes_core_sbox_inst_n1290, aes_core_sbox_inst_n1289,
         aes_core_sbox_inst_n1288, aes_core_sbox_inst_n1287,
         aes_core_sbox_inst_n1286, aes_core_sbox_inst_n1285,
         aes_core_sbox_inst_n1284, aes_core_sbox_inst_n1283,
         aes_core_sbox_inst_n1282, aes_core_sbox_inst_n1281,
         aes_core_sbox_inst_n1280, aes_core_sbox_inst_n1279,
         aes_core_sbox_inst_n1278, aes_core_sbox_inst_n1277,
         aes_core_sbox_inst_n1276, aes_core_sbox_inst_n1275,
         aes_core_sbox_inst_n1274, aes_core_sbox_inst_n1273,
         aes_core_sbox_inst_n1272, aes_core_sbox_inst_n1271,
         aes_core_sbox_inst_n1270, aes_core_sbox_inst_n1269,
         aes_core_sbox_inst_n1268, aes_core_sbox_inst_n1267,
         aes_core_sbox_inst_n1266, aes_core_sbox_inst_n1265,
         aes_core_sbox_inst_n1264, aes_core_sbox_inst_n1263,
         aes_core_sbox_inst_n1262, aes_core_sbox_inst_n1261,
         aes_core_sbox_inst_n1260, aes_core_sbox_inst_n1259,
         aes_core_sbox_inst_n1258, aes_core_sbox_inst_n1257,
         aes_core_sbox_inst_n1256, aes_core_sbox_inst_n1255,
         aes_core_sbox_inst_n1254, aes_core_sbox_inst_n1253,
         aes_core_sbox_inst_n1252, aes_core_sbox_inst_n1251,
         aes_core_sbox_inst_n1250, aes_core_sbox_inst_n1249,
         aes_core_sbox_inst_n1248, aes_core_sbox_inst_n1247,
         aes_core_sbox_inst_n1246, aes_core_sbox_inst_n1245,
         aes_core_sbox_inst_n1244, aes_core_sbox_inst_n1243,
         aes_core_sbox_inst_n1242, aes_core_sbox_inst_n1241,
         aes_core_sbox_inst_n1240, aes_core_sbox_inst_n1239,
         aes_core_sbox_inst_n1238, aes_core_sbox_inst_n1237,
         aes_core_sbox_inst_n1236, aes_core_sbox_inst_n1235,
         aes_core_sbox_inst_n1234, aes_core_sbox_inst_n1233,
         aes_core_sbox_inst_n1232, aes_core_sbox_inst_n1231,
         aes_core_sbox_inst_n1230, aes_core_sbox_inst_n1229,
         aes_core_sbox_inst_n1228, aes_core_sbox_inst_n1227,
         aes_core_sbox_inst_n1226, aes_core_sbox_inst_n1225,
         aes_core_sbox_inst_n1224, aes_core_sbox_inst_n1223,
         aes_core_sbox_inst_n1222, aes_core_sbox_inst_n1221,
         aes_core_sbox_inst_n1220, aes_core_sbox_inst_n1219,
         aes_core_sbox_inst_n1218, aes_core_sbox_inst_n1217,
         aes_core_sbox_inst_n1216, aes_core_sbox_inst_n1215,
         aes_core_sbox_inst_n1214, aes_core_sbox_inst_n1213,
         aes_core_sbox_inst_n1212, aes_core_sbox_inst_n1211,
         aes_core_sbox_inst_n1210, aes_core_sbox_inst_n1209,
         aes_core_sbox_inst_n1208, aes_core_sbox_inst_n1207,
         aes_core_sbox_inst_n1206, aes_core_sbox_inst_n1205,
         aes_core_sbox_inst_n1204, aes_core_sbox_inst_n1203,
         aes_core_sbox_inst_n1202, aes_core_sbox_inst_n1201,
         aes_core_sbox_inst_n1200, aes_core_sbox_inst_n1199,
         aes_core_sbox_inst_n1198, aes_core_sbox_inst_n1197,
         aes_core_sbox_inst_n1196, aes_core_sbox_inst_n1195,
         aes_core_sbox_inst_n1194, aes_core_sbox_inst_n1193,
         aes_core_sbox_inst_n1192, aes_core_sbox_inst_n1191,
         aes_core_sbox_inst_n1190, aes_core_sbox_inst_n1189,
         aes_core_sbox_inst_n1188, aes_core_sbox_inst_n1187,
         aes_core_sbox_inst_n1186, aes_core_sbox_inst_n1185,
         aes_core_sbox_inst_n1184, aes_core_sbox_inst_n1183,
         aes_core_sbox_inst_n1182, aes_core_sbox_inst_n1181,
         aes_core_sbox_inst_n1180, aes_core_sbox_inst_n1179,
         aes_core_sbox_inst_n1178, aes_core_sbox_inst_n1177,
         aes_core_sbox_inst_n1176, aes_core_sbox_inst_n1175,
         aes_core_sbox_inst_n1174, aes_core_sbox_inst_n1173,
         aes_core_sbox_inst_n1172, aes_core_sbox_inst_n1171,
         aes_core_sbox_inst_n1170, aes_core_sbox_inst_n1169,
         aes_core_sbox_inst_n1168, aes_core_sbox_inst_n1167,
         aes_core_sbox_inst_n1166, aes_core_sbox_inst_n1165,
         aes_core_sbox_inst_n1164, aes_core_sbox_inst_n1163,
         aes_core_sbox_inst_n1162, aes_core_sbox_inst_n1161,
         aes_core_sbox_inst_n1160, aes_core_sbox_inst_n1159,
         aes_core_sbox_inst_n1158, aes_core_sbox_inst_n1157,
         aes_core_sbox_inst_n1156, aes_core_sbox_inst_n1155,
         aes_core_sbox_inst_n1154, aes_core_sbox_inst_n1153,
         aes_core_sbox_inst_n1152, aes_core_sbox_inst_n1151,
         aes_core_sbox_inst_n1150, aes_core_sbox_inst_n1149,
         aes_core_sbox_inst_n1148, aes_core_sbox_inst_n1147,
         aes_core_sbox_inst_n1146, aes_core_sbox_inst_n1145,
         aes_core_sbox_inst_n1144, aes_core_sbox_inst_n1143,
         aes_core_sbox_inst_n1142, aes_core_sbox_inst_n1141,
         aes_core_sbox_inst_n1140, aes_core_sbox_inst_n1139,
         aes_core_sbox_inst_n1138, aes_core_sbox_inst_n1137,
         aes_core_sbox_inst_n1136, aes_core_sbox_inst_n1135,
         aes_core_sbox_inst_n1134, aes_core_sbox_inst_n1133,
         aes_core_sbox_inst_n1132, aes_core_sbox_inst_n1131,
         aes_core_sbox_inst_n1130, aes_core_sbox_inst_n1129,
         aes_core_sbox_inst_n1128, aes_core_sbox_inst_n1127,
         aes_core_sbox_inst_n1126, aes_core_sbox_inst_n1125,
         aes_core_sbox_inst_n1124, aes_core_sbox_inst_n1123,
         aes_core_sbox_inst_n1122, aes_core_sbox_inst_n1121,
         aes_core_sbox_inst_n1120, aes_core_sbox_inst_n1119,
         aes_core_sbox_inst_n1118, aes_core_sbox_inst_n1117,
         aes_core_sbox_inst_n1116, aes_core_sbox_inst_n1115,
         aes_core_sbox_inst_n1114, aes_core_sbox_inst_n1113,
         aes_core_sbox_inst_n1112, aes_core_sbox_inst_n1111,
         aes_core_sbox_inst_n1110, aes_core_sbox_inst_n1109,
         aes_core_sbox_inst_n1108, aes_core_sbox_inst_n1107,
         aes_core_sbox_inst_n1106, aes_core_sbox_inst_n1105,
         aes_core_sbox_inst_n1104, aes_core_sbox_inst_n1103,
         aes_core_sbox_inst_n1102, aes_core_sbox_inst_n1101,
         aes_core_sbox_inst_n1100, aes_core_sbox_inst_n1099,
         aes_core_sbox_inst_n1098, aes_core_sbox_inst_n1097,
         aes_core_sbox_inst_n1096, aes_core_sbox_inst_n1095,
         aes_core_sbox_inst_n1094, aes_core_sbox_inst_n1093,
         aes_core_sbox_inst_n1092, aes_core_sbox_inst_n1091,
         aes_core_sbox_inst_n1090, aes_core_sbox_inst_n1089,
         aes_core_sbox_inst_n1088, aes_core_sbox_inst_n1087,
         aes_core_sbox_inst_n1086, aes_core_sbox_inst_n1085,
         aes_core_sbox_inst_n1084, aes_core_sbox_inst_n1083,
         aes_core_sbox_inst_n1082, aes_core_sbox_inst_n1081,
         aes_core_sbox_inst_n1080, aes_core_sbox_inst_n1079,
         aes_core_sbox_inst_n1078, aes_core_sbox_inst_n1077,
         aes_core_sbox_inst_n1076, aes_core_sbox_inst_n1075,
         aes_core_sbox_inst_n1074, aes_core_sbox_inst_n1073,
         aes_core_sbox_inst_n1072, aes_core_sbox_inst_n1071,
         aes_core_sbox_inst_n1070, aes_core_sbox_inst_n1069,
         aes_core_sbox_inst_n1068, aes_core_sbox_inst_n1067,
         aes_core_sbox_inst_n1066, aes_core_sbox_inst_n1065,
         aes_core_sbox_inst_n1064, aes_core_sbox_inst_n1063,
         aes_core_sbox_inst_n1062, aes_core_sbox_inst_n1061,
         aes_core_sbox_inst_n1060, aes_core_sbox_inst_n1059,
         aes_core_sbox_inst_n1058, aes_core_sbox_inst_n1057,
         aes_core_sbox_inst_n1056, aes_core_sbox_inst_n1055,
         aes_core_sbox_inst_n1054, aes_core_sbox_inst_n1053,
         aes_core_sbox_inst_n1052, aes_core_sbox_inst_n1051,
         aes_core_sbox_inst_n1050, aes_core_sbox_inst_n1049,
         aes_core_sbox_inst_n1048, aes_core_sbox_inst_n1047,
         aes_core_sbox_inst_n1046, aes_core_sbox_inst_n1045,
         aes_core_sbox_inst_n1044, aes_core_sbox_inst_n1043,
         aes_core_sbox_inst_n1042, aes_core_sbox_inst_n1041,
         aes_core_sbox_inst_n1040, aes_core_sbox_inst_n1039,
         aes_core_sbox_inst_n1038, aes_core_sbox_inst_n1037,
         aes_core_sbox_inst_n1036, aes_core_sbox_inst_n1035,
         aes_core_sbox_inst_n1034, aes_core_sbox_inst_n1033,
         aes_core_sbox_inst_n1032, aes_core_sbox_inst_n1031,
         aes_core_sbox_inst_n1030, aes_core_sbox_inst_n1029,
         aes_core_sbox_inst_n1028, aes_core_sbox_inst_n1027,
         aes_core_sbox_inst_n1026, aes_core_sbox_inst_n1025,
         aes_core_sbox_inst_n1024, aes_core_sbox_inst_n1023,
         aes_core_sbox_inst_n1022, aes_core_sbox_inst_n1021,
         aes_core_sbox_inst_n1020, aes_core_sbox_inst_n1019,
         aes_core_sbox_inst_n1018, aes_core_sbox_inst_n1017,
         aes_core_sbox_inst_n1016, aes_core_sbox_inst_n1015,
         aes_core_sbox_inst_n1014, aes_core_sbox_inst_n1013,
         aes_core_sbox_inst_n1012, aes_core_sbox_inst_n1011,
         aes_core_sbox_inst_n1010, aes_core_sbox_inst_n1009,
         aes_core_sbox_inst_n1008, aes_core_sbox_inst_n1007,
         aes_core_sbox_inst_n1006, aes_core_sbox_inst_n1005,
         aes_core_sbox_inst_n1004, aes_core_sbox_inst_n1003,
         aes_core_sbox_inst_n1002, aes_core_sbox_inst_n1001,
         aes_core_sbox_inst_n1000, aes_core_sbox_inst_n999,
         aes_core_sbox_inst_n998, aes_core_sbox_inst_n997,
         aes_core_sbox_inst_n996, aes_core_sbox_inst_n995,
         aes_core_sbox_inst_n994, aes_core_sbox_inst_n993,
         aes_core_sbox_inst_n992, aes_core_sbox_inst_n991,
         aes_core_sbox_inst_n990, aes_core_sbox_inst_n989,
         aes_core_sbox_inst_n988, aes_core_sbox_inst_n987,
         aes_core_sbox_inst_n986, aes_core_sbox_inst_n985,
         aes_core_sbox_inst_n984, aes_core_sbox_inst_n983,
         aes_core_sbox_inst_n982, aes_core_sbox_inst_n981,
         aes_core_sbox_inst_n980, aes_core_sbox_inst_n979,
         aes_core_sbox_inst_n978, aes_core_sbox_inst_n977,
         aes_core_sbox_inst_n976, aes_core_sbox_inst_n975,
         aes_core_sbox_inst_n974, aes_core_sbox_inst_n973,
         aes_core_sbox_inst_n972, aes_core_sbox_inst_n971,
         aes_core_sbox_inst_n970, aes_core_sbox_inst_n969,
         aes_core_sbox_inst_n968, aes_core_sbox_inst_n967,
         aes_core_sbox_inst_n966, aes_core_sbox_inst_n965,
         aes_core_sbox_inst_n964, aes_core_sbox_inst_n963,
         aes_core_sbox_inst_n962, aes_core_sbox_inst_n961,
         aes_core_sbox_inst_n960, aes_core_sbox_inst_n959,
         aes_core_sbox_inst_n958, aes_core_sbox_inst_n957,
         aes_core_sbox_inst_n956, aes_core_sbox_inst_n955,
         aes_core_sbox_inst_n954, aes_core_sbox_inst_n953,
         aes_core_sbox_inst_n952, aes_core_sbox_inst_n951,
         aes_core_sbox_inst_n950, aes_core_sbox_inst_n949,
         aes_core_sbox_inst_n948, aes_core_sbox_inst_n947,
         aes_core_sbox_inst_n946, aes_core_sbox_inst_n945,
         aes_core_sbox_inst_n944, aes_core_sbox_inst_n943,
         aes_core_sbox_inst_n942, aes_core_sbox_inst_n941,
         aes_core_sbox_inst_n940, aes_core_sbox_inst_n939,
         aes_core_sbox_inst_n938, aes_core_sbox_inst_n937,
         aes_core_sbox_inst_n936, aes_core_sbox_inst_n935,
         aes_core_sbox_inst_n934, aes_core_sbox_inst_n933,
         aes_core_sbox_inst_n932, aes_core_sbox_inst_n931,
         aes_core_sbox_inst_n930, aes_core_sbox_inst_n929,
         aes_core_sbox_inst_n928, aes_core_sbox_inst_n927,
         aes_core_sbox_inst_n926, aes_core_sbox_inst_n925,
         aes_core_sbox_inst_n924, aes_core_sbox_inst_n923,
         aes_core_sbox_inst_n922, aes_core_sbox_inst_n921,
         aes_core_sbox_inst_n920, aes_core_sbox_inst_n919,
         aes_core_sbox_inst_n918, aes_core_sbox_inst_n917,
         aes_core_sbox_inst_n916, aes_core_sbox_inst_n915,
         aes_core_sbox_inst_n914, aes_core_sbox_inst_n913,
         aes_core_sbox_inst_n912, aes_core_sbox_inst_n911,
         aes_core_sbox_inst_n910, aes_core_sbox_inst_n909,
         aes_core_sbox_inst_n908, aes_core_sbox_inst_n907,
         aes_core_sbox_inst_n906, aes_core_sbox_inst_n905,
         aes_core_sbox_inst_n904, aes_core_sbox_inst_n903,
         aes_core_sbox_inst_n902, aes_core_sbox_inst_n901,
         aes_core_sbox_inst_n900, aes_core_sbox_inst_n899,
         aes_core_sbox_inst_n898, aes_core_sbox_inst_n897,
         aes_core_sbox_inst_n896, aes_core_sbox_inst_n895,
         aes_core_sbox_inst_n894, aes_core_sbox_inst_n893,
         aes_core_sbox_inst_n892, aes_core_sbox_inst_n891,
         aes_core_sbox_inst_n890, aes_core_sbox_inst_n889,
         aes_core_sbox_inst_n888, aes_core_sbox_inst_n887,
         aes_core_sbox_inst_n886, aes_core_sbox_inst_n885,
         aes_core_sbox_inst_n884, aes_core_sbox_inst_n883,
         aes_core_sbox_inst_n882, aes_core_sbox_inst_n881,
         aes_core_sbox_inst_n880, aes_core_sbox_inst_n879,
         aes_core_sbox_inst_n878, aes_core_sbox_inst_n877,
         aes_core_sbox_inst_n876, aes_core_sbox_inst_n875,
         aes_core_sbox_inst_n874, aes_core_sbox_inst_n873,
         aes_core_sbox_inst_n872, aes_core_sbox_inst_n871,
         aes_core_sbox_inst_n870, aes_core_sbox_inst_n869,
         aes_core_sbox_inst_n868, aes_core_sbox_inst_n867,
         aes_core_sbox_inst_n866, aes_core_sbox_inst_n865,
         aes_core_sbox_inst_n864, aes_core_sbox_inst_n863,
         aes_core_sbox_inst_n862, aes_core_sbox_inst_n861,
         aes_core_sbox_inst_n860, aes_core_sbox_inst_n859,
         aes_core_sbox_inst_n858, aes_core_sbox_inst_n857,
         aes_core_sbox_inst_n856, aes_core_sbox_inst_n855,
         aes_core_sbox_inst_n854, aes_core_sbox_inst_n853,
         aes_core_sbox_inst_n852, aes_core_sbox_inst_n851,
         aes_core_sbox_inst_n850, aes_core_sbox_inst_n849,
         aes_core_sbox_inst_n848, aes_core_sbox_inst_n847,
         aes_core_sbox_inst_n846, aes_core_sbox_inst_n845,
         aes_core_sbox_inst_n844, aes_core_sbox_inst_n843,
         aes_core_sbox_inst_n842, aes_core_sbox_inst_n841,
         aes_core_sbox_inst_n840, aes_core_sbox_inst_n839,
         aes_core_sbox_inst_n838, aes_core_sbox_inst_n837,
         aes_core_sbox_inst_n836, aes_core_sbox_inst_n835,
         aes_core_sbox_inst_n834, aes_core_sbox_inst_n833,
         aes_core_sbox_inst_n832, aes_core_sbox_inst_n831,
         aes_core_sbox_inst_n830, aes_core_sbox_inst_n829,
         aes_core_sbox_inst_n828, aes_core_sbox_inst_n827,
         aes_core_sbox_inst_n826, aes_core_sbox_inst_n825,
         aes_core_sbox_inst_n824, aes_core_sbox_inst_n823,
         aes_core_sbox_inst_n822, aes_core_sbox_inst_n821,
         aes_core_sbox_inst_n820, aes_core_sbox_inst_n819,
         aes_core_sbox_inst_n818, aes_core_sbox_inst_n817,
         aes_core_sbox_inst_n816, aes_core_sbox_inst_n815,
         aes_core_sbox_inst_n814, aes_core_sbox_inst_n813,
         aes_core_sbox_inst_n812, aes_core_sbox_inst_n811,
         aes_core_sbox_inst_n810, aes_core_sbox_inst_n809,
         aes_core_sbox_inst_n808, aes_core_sbox_inst_n807,
         aes_core_sbox_inst_n806, aes_core_sbox_inst_n805,
         aes_core_sbox_inst_n804, aes_core_sbox_inst_n803,
         aes_core_sbox_inst_n802, aes_core_sbox_inst_n801,
         aes_core_sbox_inst_n800, aes_core_sbox_inst_n799,
         aes_core_sbox_inst_n798, aes_core_sbox_inst_n797,
         aes_core_sbox_inst_n796, aes_core_sbox_inst_n795,
         aes_core_sbox_inst_n794, aes_core_sbox_inst_n793,
         aes_core_sbox_inst_n792, aes_core_sbox_inst_n791,
         aes_core_sbox_inst_n790, aes_core_sbox_inst_n789,
         aes_core_sbox_inst_n788, aes_core_sbox_inst_n787,
         aes_core_sbox_inst_n786, aes_core_sbox_inst_n785,
         aes_core_sbox_inst_n784, aes_core_sbox_inst_n783,
         aes_core_sbox_inst_n782, aes_core_sbox_inst_n781,
         aes_core_sbox_inst_n780, aes_core_sbox_inst_n779,
         aes_core_sbox_inst_n778, aes_core_sbox_inst_n777,
         aes_core_sbox_inst_n776, aes_core_sbox_inst_n775,
         aes_core_sbox_inst_n774, aes_core_sbox_inst_n773,
         aes_core_sbox_inst_n772, aes_core_sbox_inst_n771,
         aes_core_sbox_inst_n770, aes_core_sbox_inst_n769,
         aes_core_sbox_inst_n768, aes_core_sbox_inst_n767,
         aes_core_sbox_inst_n766, aes_core_sbox_inst_n765,
         aes_core_sbox_inst_n764, aes_core_sbox_inst_n763,
         aes_core_sbox_inst_n762, aes_core_sbox_inst_n761,
         aes_core_sbox_inst_n760, aes_core_sbox_inst_n759,
         aes_core_sbox_inst_n758, aes_core_sbox_inst_n757,
         aes_core_sbox_inst_n756, aes_core_sbox_inst_n755,
         aes_core_sbox_inst_n754, aes_core_sbox_inst_n753,
         aes_core_sbox_inst_n752, aes_core_sbox_inst_n751,
         aes_core_sbox_inst_n750, aes_core_sbox_inst_n749,
         aes_core_sbox_inst_n748, aes_core_sbox_inst_n747,
         aes_core_sbox_inst_n746, aes_core_sbox_inst_n745,
         aes_core_sbox_inst_n744, aes_core_sbox_inst_n743,
         aes_core_sbox_inst_n742, aes_core_sbox_inst_n741,
         aes_core_sbox_inst_n740, aes_core_sbox_inst_n739,
         aes_core_sbox_inst_n738, aes_core_sbox_inst_n737,
         aes_core_sbox_inst_n736, aes_core_sbox_inst_n735,
         aes_core_sbox_inst_n734, aes_core_sbox_inst_n733,
         aes_core_sbox_inst_n732, aes_core_sbox_inst_n731,
         aes_core_sbox_inst_n730, aes_core_sbox_inst_n729,
         aes_core_sbox_inst_n728, aes_core_sbox_inst_n727,
         aes_core_sbox_inst_n726, aes_core_sbox_inst_n725,
         aes_core_sbox_inst_n724, aes_core_sbox_inst_n723,
         aes_core_sbox_inst_n722, aes_core_sbox_inst_n721,
         aes_core_sbox_inst_n720, aes_core_sbox_inst_n719,
         aes_core_sbox_inst_n718, aes_core_sbox_inst_n717,
         aes_core_sbox_inst_n716, aes_core_sbox_inst_n715,
         aes_core_sbox_inst_n714, aes_core_sbox_inst_n713,
         aes_core_sbox_inst_n712, aes_core_sbox_inst_n711,
         aes_core_sbox_inst_n710, aes_core_sbox_inst_n709,
         aes_core_sbox_inst_n708, aes_core_sbox_inst_n707,
         aes_core_sbox_inst_n706, aes_core_sbox_inst_n705,
         aes_core_sbox_inst_n704, aes_core_sbox_inst_n703,
         aes_core_sbox_inst_n702, aes_core_sbox_inst_n701,
         aes_core_sbox_inst_n700, aes_core_sbox_inst_n699,
         aes_core_sbox_inst_n698, aes_core_sbox_inst_n697,
         aes_core_sbox_inst_n696, aes_core_sbox_inst_n695,
         aes_core_sbox_inst_n694, aes_core_sbox_inst_n693,
         aes_core_sbox_inst_n692, aes_core_sbox_inst_n691,
         aes_core_sbox_inst_n690, aes_core_sbox_inst_n689,
         aes_core_sbox_inst_n688, aes_core_sbox_inst_n687,
         aes_core_sbox_inst_n686, aes_core_sbox_inst_n685,
         aes_core_sbox_inst_n684, aes_core_sbox_inst_n683,
         aes_core_sbox_inst_n682, aes_core_sbox_inst_n681,
         aes_core_sbox_inst_n680, aes_core_sbox_inst_n679,
         aes_core_sbox_inst_n678, aes_core_sbox_inst_n677,
         aes_core_sbox_inst_n676, aes_core_sbox_inst_n675,
         aes_core_sbox_inst_n674, aes_core_sbox_inst_n673,
         aes_core_sbox_inst_n672, aes_core_sbox_inst_n671,
         aes_core_sbox_inst_n670, aes_core_sbox_inst_n669,
         aes_core_sbox_inst_n668, aes_core_sbox_inst_n667,
         aes_core_sbox_inst_n666, aes_core_sbox_inst_n665,
         aes_core_sbox_inst_n664, aes_core_sbox_inst_n663,
         aes_core_sbox_inst_n662, aes_core_sbox_inst_n661,
         aes_core_sbox_inst_n660, aes_core_sbox_inst_n659,
         aes_core_sbox_inst_n658, aes_core_sbox_inst_n657,
         aes_core_sbox_inst_n656, aes_core_sbox_inst_n655,
         aes_core_sbox_inst_n654, aes_core_sbox_inst_n653,
         aes_core_sbox_inst_n652, aes_core_sbox_inst_n651,
         aes_core_sbox_inst_n650, aes_core_sbox_inst_n649,
         aes_core_sbox_inst_n648, aes_core_sbox_inst_n647,
         aes_core_sbox_inst_n646, aes_core_sbox_inst_n645,
         aes_core_sbox_inst_n644, aes_core_sbox_inst_n643,
         aes_core_sbox_inst_n642, aes_core_sbox_inst_n641,
         aes_core_sbox_inst_n640, aes_core_sbox_inst_n639,
         aes_core_sbox_inst_n638, aes_core_sbox_inst_n637,
         aes_core_sbox_inst_n636, aes_core_sbox_inst_n635,
         aes_core_sbox_inst_n634, aes_core_sbox_inst_n633,
         aes_core_sbox_inst_n632, aes_core_sbox_inst_n631,
         aes_core_sbox_inst_n630, aes_core_sbox_inst_n629,
         aes_core_sbox_inst_n628, aes_core_sbox_inst_n627,
         aes_core_sbox_inst_n626, aes_core_sbox_inst_n625,
         aes_core_sbox_inst_n624, aes_core_sbox_inst_n623,
         aes_core_sbox_inst_n622, aes_core_sbox_inst_n621,
         aes_core_sbox_inst_n620, aes_core_sbox_inst_n619,
         aes_core_sbox_inst_n618, aes_core_sbox_inst_n616,
         aes_core_sbox_inst_n615, aes_core_sbox_inst_n614,
         aes_core_sbox_inst_n613, aes_core_sbox_inst_n612,
         aes_core_sbox_inst_n611, aes_core_sbox_inst_n610,
         aes_core_sbox_inst_n609, aes_core_sbox_inst_n608,
         aes_core_sbox_inst_n607, aes_core_sbox_inst_n606,
         aes_core_sbox_inst_n605, aes_core_sbox_inst_n604,
         aes_core_sbox_inst_n603, aes_core_sbox_inst_n602,
         aes_core_sbox_inst_n601, aes_core_sbox_inst_n600,
         aes_core_sbox_inst_n599, aes_core_sbox_inst_n598,
         aes_core_sbox_inst_n597, aes_core_sbox_inst_n596,
         aes_core_sbox_inst_n595, aes_core_sbox_inst_n594,
         aes_core_sbox_inst_n593, aes_core_sbox_inst_n592,
         aes_core_sbox_inst_n591, aes_core_sbox_inst_n590,
         aes_core_sbox_inst_n589, aes_core_sbox_inst_n588,
         aes_core_sbox_inst_n587, aes_core_sbox_inst_n586,
         aes_core_sbox_inst_n585, aes_core_sbox_inst_n584,
         aes_core_sbox_inst_n583, aes_core_sbox_inst_n582,
         aes_core_sbox_inst_n581, aes_core_sbox_inst_n580,
         aes_core_sbox_inst_n579, aes_core_sbox_inst_n578,
         aes_core_sbox_inst_n577, aes_core_sbox_inst_n576,
         aes_core_sbox_inst_n575, aes_core_sbox_inst_n574,
         aes_core_sbox_inst_n573, aes_core_sbox_inst_n572,
         aes_core_sbox_inst_n571, aes_core_sbox_inst_n570,
         aes_core_sbox_inst_n569, aes_core_sbox_inst_n568,
         aes_core_sbox_inst_n567, aes_core_sbox_inst_n566,
         aes_core_sbox_inst_n565, aes_core_sbox_inst_n564,
         aes_core_sbox_inst_n563, aes_core_sbox_inst_n562,
         aes_core_sbox_inst_n561, aes_core_sbox_inst_n560,
         aes_core_sbox_inst_n559, aes_core_sbox_inst_n558,
         aes_core_sbox_inst_n557, aes_core_sbox_inst_n556,
         aes_core_sbox_inst_n555, aes_core_sbox_inst_n554,
         aes_core_sbox_inst_n553, aes_core_sbox_inst_n552,
         aes_core_sbox_inst_n551, aes_core_sbox_inst_n550,
         aes_core_sbox_inst_n549, aes_core_sbox_inst_n548,
         aes_core_sbox_inst_n547, aes_core_sbox_inst_n546,
         aes_core_sbox_inst_n545, aes_core_sbox_inst_n544,
         aes_core_sbox_inst_n543, aes_core_sbox_inst_n542,
         aes_core_sbox_inst_n541, aes_core_sbox_inst_n540,
         aes_core_sbox_inst_n539, aes_core_sbox_inst_n538,
         aes_core_sbox_inst_n537, aes_core_sbox_inst_n536,
         aes_core_sbox_inst_n535, aes_core_sbox_inst_n534,
         aes_core_sbox_inst_n533, aes_core_sbox_inst_n532,
         aes_core_sbox_inst_n531, aes_core_sbox_inst_n530,
         aes_core_sbox_inst_n529, aes_core_sbox_inst_n528,
         aes_core_sbox_inst_n527, aes_core_sbox_inst_n526,
         aes_core_sbox_inst_n525, aes_core_sbox_inst_n524,
         aes_core_sbox_inst_n523, aes_core_sbox_inst_n522,
         aes_core_sbox_inst_n521, aes_core_sbox_inst_n520,
         aes_core_sbox_inst_n519, aes_core_sbox_inst_n518,
         aes_core_sbox_inst_n517, aes_core_sbox_inst_n516,
         aes_core_sbox_inst_n515, aes_core_sbox_inst_n514,
         aes_core_sbox_inst_n513, aes_core_sbox_inst_n512,
         aes_core_sbox_inst_n511, aes_core_sbox_inst_n510,
         aes_core_sbox_inst_n509, aes_core_sbox_inst_n508,
         aes_core_sbox_inst_n507, aes_core_sbox_inst_n506,
         aes_core_sbox_inst_n505, aes_core_sbox_inst_n504,
         aes_core_sbox_inst_n503, aes_core_sbox_inst_n502,
         aes_core_sbox_inst_n501, aes_core_sbox_inst_n500,
         aes_core_sbox_inst_n499, aes_core_sbox_inst_n498,
         aes_core_sbox_inst_n497, aes_core_sbox_inst_n496,
         aes_core_sbox_inst_n495, aes_core_sbox_inst_n494,
         aes_core_sbox_inst_n493, aes_core_sbox_inst_n492,
         aes_core_sbox_inst_n491, aes_core_sbox_inst_n490,
         aes_core_sbox_inst_n489, aes_core_sbox_inst_n488,
         aes_core_sbox_inst_n487, aes_core_sbox_inst_n486,
         aes_core_sbox_inst_n485, aes_core_sbox_inst_n484,
         aes_core_sbox_inst_n483, aes_core_sbox_inst_n482,
         aes_core_sbox_inst_n481, aes_core_sbox_inst_n480,
         aes_core_sbox_inst_n479, aes_core_sbox_inst_n478,
         aes_core_sbox_inst_n477, aes_core_sbox_inst_n476,
         aes_core_sbox_inst_n475, aes_core_sbox_inst_n474,
         aes_core_sbox_inst_n473, aes_core_sbox_inst_n472,
         aes_core_sbox_inst_n471, aes_core_sbox_inst_n470,
         aes_core_sbox_inst_n469, aes_core_sbox_inst_n468,
         aes_core_sbox_inst_n467, aes_core_sbox_inst_n466,
         aes_core_sbox_inst_n465, aes_core_sbox_inst_n464,
         aes_core_sbox_inst_n463, aes_core_sbox_inst_n462,
         aes_core_sbox_inst_n461, aes_core_sbox_inst_n460,
         aes_core_sbox_inst_n459, aes_core_sbox_inst_n458,
         aes_core_sbox_inst_n457, aes_core_sbox_inst_n456,
         aes_core_sbox_inst_n455, aes_core_sbox_inst_n454,
         aes_core_sbox_inst_n453, aes_core_sbox_inst_n452,
         aes_core_sbox_inst_n451, aes_core_sbox_inst_n449,
         aes_core_sbox_inst_n448, aes_core_sbox_inst_n447,
         aes_core_sbox_inst_n446, aes_core_sbox_inst_n445,
         aes_core_sbox_inst_n444, aes_core_sbox_inst_n443,
         aes_core_sbox_inst_n442, aes_core_sbox_inst_n441,
         aes_core_sbox_inst_n440, aes_core_sbox_inst_n439,
         aes_core_sbox_inst_n438, aes_core_sbox_inst_n437,
         aes_core_sbox_inst_n436, aes_core_sbox_inst_n435,
         aes_core_sbox_inst_n434, aes_core_sbox_inst_n433,
         aes_core_sbox_inst_n432, aes_core_sbox_inst_n431,
         aes_core_sbox_inst_n430, aes_core_sbox_inst_n429,
         aes_core_sbox_inst_n428, aes_core_sbox_inst_n427,
         aes_core_sbox_inst_n426, aes_core_sbox_inst_n425,
         aes_core_sbox_inst_n424, aes_core_sbox_inst_n423,
         aes_core_sbox_inst_n422, aes_core_sbox_inst_n421,
         aes_core_sbox_inst_n420, aes_core_sbox_inst_n419,
         aes_core_sbox_inst_n418, aes_core_sbox_inst_n417,
         aes_core_sbox_inst_n416, aes_core_sbox_inst_n415,
         aes_core_sbox_inst_n414, aes_core_sbox_inst_n413,
         aes_core_sbox_inst_n412, aes_core_sbox_inst_n411,
         aes_core_sbox_inst_n410, aes_core_sbox_inst_n409,
         aes_core_sbox_inst_n408, aes_core_sbox_inst_n407,
         aes_core_sbox_inst_n406, aes_core_sbox_inst_n405,
         aes_core_sbox_inst_n404, aes_core_sbox_inst_n403,
         aes_core_sbox_inst_n402, aes_core_sbox_inst_n401,
         aes_core_sbox_inst_n400, aes_core_sbox_inst_n399,
         aes_core_sbox_inst_n398, aes_core_sbox_inst_n397,
         aes_core_sbox_inst_n396, aes_core_sbox_inst_n395,
         aes_core_sbox_inst_n394, aes_core_sbox_inst_n393,
         aes_core_sbox_inst_n392, aes_core_sbox_inst_n391,
         aes_core_sbox_inst_n390, aes_core_sbox_inst_n389,
         aes_core_sbox_inst_n388, aes_core_sbox_inst_n387,
         aes_core_sbox_inst_n386, aes_core_sbox_inst_n385,
         aes_core_sbox_inst_n384, aes_core_sbox_inst_n383,
         aes_core_sbox_inst_n382, aes_core_sbox_inst_n381,
         aes_core_sbox_inst_n380, aes_core_sbox_inst_n379,
         aes_core_sbox_inst_n378, aes_core_sbox_inst_n377,
         aes_core_sbox_inst_n376, aes_core_sbox_inst_n375,
         aes_core_sbox_inst_n374, aes_core_sbox_inst_n373,
         aes_core_sbox_inst_n372, aes_core_sbox_inst_n371,
         aes_core_sbox_inst_n370, aes_core_sbox_inst_n369,
         aes_core_sbox_inst_n368, aes_core_sbox_inst_n367,
         aes_core_sbox_inst_n366, aes_core_sbox_inst_n365,
         aes_core_sbox_inst_n364, aes_core_sbox_inst_n363,
         aes_core_sbox_inst_n362, aes_core_sbox_inst_n361,
         aes_core_sbox_inst_n360, aes_core_sbox_inst_n359,
         aes_core_sbox_inst_n358, aes_core_sbox_inst_n357,
         aes_core_sbox_inst_n356, aes_core_sbox_inst_n355,
         aes_core_sbox_inst_n354, aes_core_sbox_inst_n353,
         aes_core_sbox_inst_n352, aes_core_sbox_inst_n351,
         aes_core_sbox_inst_n350, aes_core_sbox_inst_n349,
         aes_core_sbox_inst_n348, aes_core_sbox_inst_n347,
         aes_core_sbox_inst_n346, aes_core_sbox_inst_n345,
         aes_core_sbox_inst_n344, aes_core_sbox_inst_n343,
         aes_core_sbox_inst_n342, aes_core_sbox_inst_n341,
         aes_core_sbox_inst_n340, aes_core_sbox_inst_n339,
         aes_core_sbox_inst_n338, aes_core_sbox_inst_n337,
         aes_core_sbox_inst_n336, aes_core_sbox_inst_n335,
         aes_core_sbox_inst_n334, aes_core_sbox_inst_n333,
         aes_core_sbox_inst_n332, aes_core_sbox_inst_n331,
         aes_core_sbox_inst_n330, aes_core_sbox_inst_n329,
         aes_core_sbox_inst_n328, aes_core_sbox_inst_n327,
         aes_core_sbox_inst_n326, aes_core_sbox_inst_n325,
         aes_core_sbox_inst_n324, aes_core_sbox_inst_n323,
         aes_core_sbox_inst_n322, aes_core_sbox_inst_n321,
         aes_core_sbox_inst_n320, aes_core_sbox_inst_n319,
         aes_core_sbox_inst_n318, aes_core_sbox_inst_n317,
         aes_core_sbox_inst_n315, aes_core_sbox_inst_n314,
         aes_core_sbox_inst_n313, aes_core_sbox_inst_n312,
         aes_core_sbox_inst_n311, aes_core_sbox_inst_n310,
         aes_core_sbox_inst_n309, aes_core_sbox_inst_n308,
         aes_core_sbox_inst_n307, aes_core_sbox_inst_n306,
         aes_core_sbox_inst_n305, aes_core_sbox_inst_n304,
         aes_core_sbox_inst_n303, aes_core_sbox_inst_n302,
         aes_core_sbox_inst_n301, aes_core_sbox_inst_n300,
         aes_core_sbox_inst_n299, aes_core_sbox_inst_n298,
         aes_core_sbox_inst_n297, aes_core_sbox_inst_n296,
         aes_core_sbox_inst_n295, aes_core_sbox_inst_n294,
         aes_core_sbox_inst_n293, aes_core_sbox_inst_n292,
         aes_core_sbox_inst_n291, aes_core_sbox_inst_n290,
         aes_core_sbox_inst_n289, aes_core_sbox_inst_n288,
         aes_core_sbox_inst_n287, aes_core_sbox_inst_n286,
         aes_core_sbox_inst_n285, aes_core_sbox_inst_n284,
         aes_core_sbox_inst_n283, aes_core_sbox_inst_n282,
         aes_core_sbox_inst_n281, aes_core_sbox_inst_n280,
         aes_core_sbox_inst_n279, aes_core_sbox_inst_n278,
         aes_core_sbox_inst_n277, aes_core_sbox_inst_n276,
         aes_core_sbox_inst_n275, aes_core_sbox_inst_n274,
         aes_core_sbox_inst_n272, aes_core_sbox_inst_n271,
         aes_core_sbox_inst_n270, aes_core_sbox_inst_n269,
         aes_core_sbox_inst_n268, aes_core_sbox_inst_n267,
         aes_core_sbox_inst_n266, aes_core_sbox_inst_n265,
         aes_core_sbox_inst_n264, aes_core_sbox_inst_n263,
         aes_core_sbox_inst_n262, aes_core_sbox_inst_n261,
         aes_core_sbox_inst_n260, reg_in_n1032, reg_in_n1031, reg_in_n1030,
         reg_in_n1029, reg_in_n1028, reg_in_n1027, reg_in_n1026, reg_in_n1025,
         reg_in_n1024, reg_in_n1023, reg_in_n1022, reg_in_n1021, reg_in_n1020,
         reg_in_n1019, reg_in_n1018, reg_in_n1017, reg_in_n1016, reg_in_n1015,
         reg_in_n1014, reg_in_n1013, reg_in_n1012, reg_in_n1011, reg_in_n1010,
         reg_in_n1009, reg_in_n1008, reg_in_n1007, reg_in_n1006, reg_in_n1005,
         reg_in_n1004, reg_in_n1003, reg_in_n1002, reg_in_n1001, reg_in_n1000,
         reg_in_n999, reg_in_n998, reg_in_n997, reg_in_n996, reg_in_n995,
         reg_in_n994, reg_in_n993, reg_in_n992, reg_in_n991, reg_in_n990,
         reg_in_n989, reg_in_n988, reg_in_n987, reg_in_n986, reg_in_n985,
         reg_in_n984, reg_in_n983, reg_in_n982, reg_in_n981, reg_in_n980,
         reg_in_n979, reg_in_n978, reg_in_n977, reg_in_n976, reg_in_n975,
         reg_in_n974, reg_in_n973, reg_in_n972, reg_in_n971, reg_in_n970,
         reg_in_n969, reg_in_n968, reg_in_n967, reg_in_n966, reg_in_n965,
         reg_in_n964, reg_in_n963, reg_in_n962, reg_in_n961, reg_in_n960,
         reg_in_n959, reg_in_n958, reg_in_n957, reg_in_n956, reg_in_n955,
         reg_in_n954, reg_in_n953, reg_in_n952, reg_in_n951, reg_in_n950,
         reg_in_n949, reg_in_n948, reg_in_n947, reg_in_n946, reg_in_n945,
         reg_in_n944, reg_in_n943, reg_in_n942, reg_in_n941, reg_in_n940,
         reg_in_n939, reg_in_n938, reg_in_n937, reg_in_n936, reg_in_n935,
         reg_in_n934, reg_in_n933, reg_in_n932, reg_in_n931, reg_in_n930,
         reg_in_n929, reg_in_n928, reg_in_n927, reg_in_n926, reg_in_n925,
         reg_in_n924, reg_in_n923, reg_in_n922, reg_in_n921, reg_in_n920,
         reg_in_n919, reg_in_n918, reg_in_n917, reg_in_n916, reg_in_n915,
         reg_in_n914, reg_in_n913, reg_in_n912, reg_in_n911, reg_in_n910,
         reg_in_n909, reg_in_n908, reg_in_n907, reg_in_n906, reg_in_n905,
         reg_in_n904, reg_in_n903, reg_in_n902, reg_in_n901, reg_in_n900,
         reg_in_n899, reg_in_n898, reg_in_n897, reg_in_n896, reg_in_n895,
         reg_in_n894, reg_in_n893, reg_in_n892, reg_in_n891, reg_in_n890,
         reg_in_n889, reg_in_n888, reg_in_n887, reg_in_n886, reg_in_n885,
         reg_in_n884, reg_in_n883, reg_in_n882, reg_in_n881, reg_in_n880,
         reg_in_n879, reg_in_n878, reg_in_n877, reg_in_n876, reg_in_n875,
         reg_in_n874, reg_in_n873, reg_in_n872, reg_in_n871, reg_in_n870,
         reg_in_n869, reg_in_n868, reg_in_n867, reg_in_n866, reg_in_n865,
         reg_in_n864, reg_in_n863, reg_in_n862, reg_in_n861, reg_in_n860,
         reg_in_n859, reg_in_n858, reg_in_n857, reg_in_n856, reg_in_n855,
         reg_in_n854, reg_in_n853, reg_in_n852, reg_in_n851, reg_in_n850,
         reg_in_n849, reg_in_n848, reg_in_n847, reg_in_n846, reg_in_n845,
         reg_in_n844, reg_in_n843, reg_in_n842, reg_in_n841, reg_in_n840,
         reg_in_n839, reg_in_n838, reg_in_n837, reg_in_n836, reg_in_n835,
         reg_in_n834, reg_in_n833, reg_in_n832, reg_in_n831, reg_in_n830,
         reg_in_n829, reg_in_n828, reg_in_n827, reg_in_n826, reg_in_n825,
         reg_in_n824, reg_in_n823, reg_in_n822, reg_in_n821, reg_in_n820,
         reg_in_n819, reg_in_n818, reg_in_n817, reg_in_n816, reg_in_n815,
         reg_in_n814, reg_in_n813, reg_in_n812, reg_in_n811, reg_in_n810,
         reg_in_n809, reg_in_n808, reg_in_n807, reg_in_n806, reg_in_n805,
         reg_in_n804, reg_in_n803, reg_in_n802, reg_in_n801, reg_in_n800,
         reg_in_n799, reg_in_n798, reg_in_n797, reg_in_n796, reg_in_n795,
         reg_in_n794, reg_in_n793, reg_in_n792, reg_in_n791, reg_in_n790,
         reg_in_n789, reg_in_n788, reg_in_n787, reg_in_n786, reg_in_n785,
         reg_in_n784, reg_in_n783, reg_in_n782, reg_in_n781, reg_in_n780,
         reg_in_n779, reg_in_n778, reg_in_n777, reg_in_n776, reg_in_n775,
         reg_in_n774, reg_in_n773, reg_in_n772, reg_in_n259, reg_in_n257,
         reg_in_n256, reg_in_n255, reg_in_n254, reg_in_n253, reg_in_n252,
         reg_in_n251, reg_in_n250, reg_in_n249, reg_in_n248, reg_in_n247,
         reg_in_n246, reg_in_n245, reg_in_n244, reg_in_n243, reg_in_n242,
         reg_in_n241, reg_in_n240, reg_in_n239, reg_in_n238, reg_in_n237,
         reg_in_n236, reg_in_n235, reg_in_n234, reg_in_n233, reg_in_n232,
         reg_in_n231, reg_in_n230, reg_in_n229, reg_in_n228, reg_in_n227,
         reg_in_n226, reg_in_n225, reg_in_n224, reg_in_n223, reg_in_n222,
         reg_in_n221, reg_in_n220, reg_in_n219, reg_in_n218, reg_in_n217,
         reg_in_n216, reg_in_n215, reg_in_n214, reg_in_n213, reg_in_n212,
         reg_in_n211, reg_in_n210, reg_in_n209, reg_in_n208, reg_in_n207,
         reg_in_n206, reg_in_n205, reg_in_n204, reg_in_n203, reg_in_n202,
         reg_in_n201, reg_in_n200, reg_in_n199, reg_in_n198, reg_in_n197,
         reg_in_n196, reg_in_n195, reg_in_n194, reg_in_n193, reg_in_n192,
         reg_in_n191, reg_in_n190, reg_in_n189, reg_in_n188, reg_in_n187,
         reg_in_n186, reg_in_n185, reg_in_n184, reg_in_n183, reg_in_n182,
         reg_in_n181, reg_in_n180, reg_in_n179, reg_in_n178, reg_in_n177,
         reg_in_n176, reg_in_n175, reg_in_n174, reg_in_n173, reg_in_n172,
         reg_in_n171, reg_in_n170, reg_in_n169, reg_in_n168, reg_in_n167,
         reg_in_n166, reg_in_n165, reg_in_n164, reg_in_n163, reg_in_n162,
         reg_in_n161, reg_in_n160, reg_in_n159, reg_in_n158, reg_in_n157,
         reg_in_n156, reg_in_n155, reg_in_n154, reg_in_n153, reg_in_n152,
         reg_in_n151, reg_in_n150, reg_in_n149, reg_in_n148, reg_in_n147,
         reg_in_n146, reg_in_n145, reg_in_n144, reg_in_n143, reg_in_n142,
         reg_in_n141, reg_in_n140, reg_in_n139, reg_in_n138, reg_in_n137,
         reg_in_n136, reg_in_n135, reg_in_n134, reg_in_n133, reg_in_n132,
         reg_in_n131, reg_in_n130, reg_in_n129, reg_in_n128, reg_in_n127,
         reg_in_n126, reg_in_n125, reg_in_n124, reg_in_n123, reg_in_n122,
         reg_in_n121, reg_in_n120, reg_in_n119, reg_in_n118, reg_in_n117,
         reg_in_n116, reg_in_n115, reg_in_n114, reg_in_n113, reg_in_n112,
         reg_in_n111, reg_in_n110, reg_in_n109, reg_in_n108, reg_in_n107,
         reg_in_n106, reg_in_n105, reg_in_n104, reg_in_n103, reg_in_n102,
         reg_in_n101, reg_in_n100, reg_in_n99, reg_in_n98, reg_in_n97,
         reg_in_n96, reg_in_n95, reg_in_n94, reg_in_n93, reg_in_n92,
         reg_in_n91, reg_in_n90, reg_in_n89, reg_in_n88, reg_in_n87,
         reg_in_n86, reg_in_n85, reg_in_n84, reg_in_n83, reg_in_n82,
         reg_in_n81, reg_in_n80, reg_in_n79, reg_in_n78, reg_in_n77,
         reg_in_n76, reg_in_n75, reg_in_n74, reg_in_n73, reg_in_n72,
         reg_in_n71, reg_in_n70, reg_in_n69, reg_in_n68, reg_in_n67,
         reg_in_n66, reg_in_n65, reg_in_n64, reg_in_n63, reg_in_n62,
         reg_in_n61, reg_in_n60, reg_in_n59, reg_in_n58, reg_in_n57,
         reg_in_n56, reg_in_n55, reg_in_n54, reg_in_n53, reg_in_n52,
         reg_in_n51, reg_in_n50, reg_in_n49, reg_in_n48, reg_in_n47,
         reg_in_n46, reg_in_n45, reg_in_n44, reg_in_n43, reg_in_n42,
         reg_in_n41, reg_in_n40, reg_in_n39, reg_in_n38, reg_in_n37,
         reg_in_n36, reg_in_n35, reg_in_n34, reg_in_n33, reg_in_n32,
         reg_in_n31, reg_in_n30, reg_in_n29, reg_in_n28, reg_in_n27,
         reg_in_n26, reg_in_n25, reg_in_n24, reg_in_n23, reg_in_n22,
         reg_in_n21, reg_in_n20, reg_in_n19, reg_in_n18, reg_in_n17,
         reg_in_n16, reg_in_n15, reg_in_n14, reg_in_n13, reg_in_n12,
         reg_in_n11, reg_in_n10, reg_in_n9, reg_in_n8, reg_in_n7, reg_in_n6,
         reg_in_n5, reg_in_n4, reg_in_n3, reg_in_n2, reg_in_n771, reg_in_n770,
         reg_in_n769, reg_in_n768, reg_in_n767, reg_in_n766, reg_in_n765,
         reg_in_n764, reg_in_n763, reg_in_n762, reg_in_n761, reg_in_n760,
         reg_in_n759, reg_in_n758, reg_in_n757, reg_in_n756, reg_in_n755,
         reg_in_n754, reg_in_n753, reg_in_n752, reg_in_n751, reg_in_n750,
         reg_in_n749, reg_in_n748, reg_in_n747, reg_in_n746, reg_in_n745,
         reg_in_n744, reg_in_n743, reg_in_n742, reg_in_n741, reg_in_n740,
         reg_in_n739, reg_in_n738, reg_in_n737, reg_in_n736, reg_in_n735,
         reg_in_n734, reg_in_n733, reg_in_n732, reg_in_n731, reg_in_n730,
         reg_in_n729, reg_in_n728, reg_in_n727, reg_in_n726, reg_in_n725,
         reg_in_n724, reg_in_n723, reg_in_n722, reg_in_n721, reg_in_n720,
         reg_in_n719, reg_in_n718, reg_in_n717, reg_in_n716, reg_in_n715,
         reg_in_n714, reg_in_n713, reg_in_n712, reg_in_n711, reg_in_n710,
         reg_in_n709, reg_in_n708, reg_in_n707, reg_in_n706, reg_in_n705,
         reg_in_n704, reg_in_n703, reg_in_n702, reg_in_n701, reg_in_n700,
         reg_in_n699, reg_in_n698, reg_in_n697, reg_in_n696, reg_in_n695,
         reg_in_n694, reg_in_n693, reg_in_n692, reg_in_n691, reg_in_n690,
         reg_in_n689, reg_in_n688, reg_in_n687, reg_in_n686, reg_in_n685,
         reg_in_n684, reg_in_n683, reg_in_n682, reg_in_n681, reg_in_n680,
         reg_in_n679, reg_in_n678, reg_in_n677, reg_in_n676, reg_in_n675,
         reg_in_n674, reg_in_n673, reg_in_n672, reg_in_n671, reg_in_n670,
         reg_in_n669, reg_in_n668, reg_in_n667, reg_in_n666, reg_in_n665,
         reg_in_n664, reg_in_n663, reg_in_n662, reg_in_n661, reg_in_n660,
         reg_in_n659, reg_in_n658, reg_in_n657, reg_in_n656, reg_in_n655,
         reg_in_n654, reg_in_n653, reg_in_n652, reg_in_n651, reg_in_n650,
         reg_in_n649, reg_in_n648, reg_in_n647, reg_in_n646, reg_in_n645,
         reg_in_n644, reg_in_n643, reg_in_n642, reg_in_n641, reg_in_n640,
         reg_in_n639, reg_in_n638, reg_in_n637, reg_in_n636, reg_in_n635,
         reg_in_n634, reg_in_n633, reg_in_n632, reg_in_n631, reg_in_n630,
         reg_in_n629, reg_in_n628, reg_in_n627, reg_in_n626, reg_in_n625,
         reg_in_n624, reg_in_n623, reg_in_n622, reg_in_n621, reg_in_n620,
         reg_in_n619, reg_in_n618, reg_in_n617, reg_in_n616, reg_in_n615,
         reg_in_n614, reg_in_n613, reg_in_n612, reg_in_n611, reg_in_n610,
         reg_in_n609, reg_in_n608, reg_in_n607, reg_in_n606, reg_in_n605,
         reg_in_n604, reg_in_n603, reg_in_n602, reg_in_n601, reg_in_n600,
         reg_in_n599, reg_in_n598, reg_in_n597, reg_in_n596, reg_in_n595,
         reg_in_n594, reg_in_n593, reg_in_n592, reg_in_n591, reg_in_n590,
         reg_in_n589, reg_in_n588, reg_in_n587, reg_in_n586, reg_in_n585,
         reg_in_n584, reg_in_n583, reg_in_n582, reg_in_n581, reg_in_n580,
         reg_in_n579, reg_in_n578, reg_in_n577, reg_in_n576, reg_in_n575,
         reg_in_n574, reg_in_n573, reg_in_n572, reg_in_n571, reg_in_n570,
         reg_in_n569, reg_in_n568, reg_in_n567, reg_in_n566, reg_in_n565,
         reg_in_n564, reg_in_n563, reg_in_n562, reg_in_n561, reg_in_n560,
         reg_in_n559, reg_in_n558, reg_in_n557, reg_in_n556, reg_in_n555,
         reg_in_n554, reg_in_n553, reg_in_n552, reg_in_n551, reg_in_n550,
         reg_in_n549, reg_in_n548, reg_in_n547, reg_in_n546, reg_in_n545,
         reg_in_n544, reg_in_n543, reg_in_n542, reg_in_n541, reg_in_n540,
         reg_in_n539, reg_in_n538, reg_in_n537, reg_in_n536, reg_in_n535,
         reg_in_n534, reg_in_n533, reg_in_n532, reg_in_n531, reg_in_n530,
         reg_in_n529, reg_in_n528, reg_in_n527, reg_in_n526, reg_in_n525,
         reg_in_n524, reg_in_n523, reg_in_n522, reg_in_n521, reg_in_n520,
         reg_in_n519, reg_in_n518, reg_in_n517, reg_in_n516, reg_in_n515,
         reg_in_n514, reg_in_n513, reg_in_n512, reg_in_n511, reg_in_n510,
         reg_in_n509, reg_in_n508, reg_in_n507, reg_in_n506, reg_in_n505,
         reg_in_n504, reg_in_n503, reg_in_n502, reg_in_n501, reg_in_n500,
         reg_in_n499, reg_in_n498, reg_in_n497, reg_in_n496, reg_in_n495,
         reg_in_n494, reg_in_n493, reg_in_n492, reg_in_n491, reg_in_n490,
         reg_in_n489, reg_in_n488, reg_in_n487, reg_in_n486, reg_in_n485,
         reg_in_n484, reg_in_n483, reg_in_n482, reg_in_n481, reg_in_n480,
         reg_in_n479, reg_in_n478, reg_in_n477, reg_in_n476, reg_in_n475,
         reg_in_n474, reg_in_n473, reg_in_n472, reg_in_n471, reg_in_n470,
         reg_in_n469, reg_in_n468, reg_in_n467, reg_in_n466, reg_in_n465,
         reg_in_n464, reg_in_n463, reg_in_n462, reg_in_n461, reg_in_n460,
         reg_in_n459, reg_in_n458, reg_in_n457, reg_in_n456, reg_in_n455,
         reg_in_n454, reg_in_n453, reg_in_n452, reg_in_n451, reg_in_n450,
         reg_in_n449, reg_in_n448, reg_in_n447, reg_in_n446, reg_in_n445,
         reg_in_n444, reg_in_n443, reg_in_n442, reg_in_n441, reg_in_n440,
         reg_in_n439, reg_in_n438, reg_in_n437, reg_in_n436, reg_in_n435,
         reg_in_n434, reg_in_n433, reg_in_n432, reg_in_n431, reg_in_n430,
         reg_in_n429, reg_in_n428, reg_in_n427, reg_in_n426, reg_in_n425,
         reg_in_n424, reg_in_n423, reg_in_n422, reg_in_n421, reg_in_n420,
         reg_in_n419, reg_in_n418, reg_in_n417, reg_in_n416, reg_in_n415,
         reg_in_n414, reg_in_n413, reg_in_n412, reg_in_n411, reg_in_n410,
         reg_in_n409, reg_in_n408, reg_in_n407, reg_in_n406, reg_in_n405,
         reg_in_n404, reg_in_n403, reg_in_n402, reg_in_n401, reg_in_n400,
         reg_in_n399, reg_in_n398, reg_in_n397, reg_in_n396, reg_in_n395,
         reg_in_n394, reg_in_n393, reg_in_n392, reg_in_n391, reg_in_n390,
         reg_in_n389, reg_in_n388, reg_in_n387, reg_in_n386, reg_in_n385,
         reg_in_n384, reg_in_n383, reg_in_n382, reg_in_n381, reg_in_n380,
         reg_in_n379, reg_in_n378, reg_in_n377, reg_in_n376, reg_in_n375,
         reg_in_n374, reg_in_n373, reg_in_n372, reg_in_n371, reg_in_n370,
         reg_in_n369, reg_in_n368, reg_in_n367, reg_in_n366, reg_in_n365,
         reg_in_n364, reg_in_n363, reg_in_n362, reg_in_n361, reg_in_n360,
         reg_in_n359, reg_in_n358, reg_in_n357, reg_in_n356, reg_in_n355,
         reg_in_n354, reg_in_n353, reg_in_n352, reg_in_n351, reg_in_n350,
         reg_in_n349, reg_in_n348, reg_in_n347, reg_in_n346, reg_in_n345,
         reg_in_n344, reg_in_n343, reg_in_n342, reg_in_n341, reg_in_n340,
         reg_in_n339, reg_in_n338, reg_in_n337, reg_in_n336, reg_in_n335,
         reg_in_n334, reg_in_n333, reg_in_n332, reg_in_n331, reg_in_n330,
         reg_in_n329, reg_in_n328, reg_in_n327, reg_in_n326, reg_in_n325,
         reg_in_n324, reg_in_n323, reg_in_n322, reg_in_n321, reg_in_n320,
         reg_in_n319, reg_in_n318, reg_in_n317, reg_in_n316, reg_in_n315,
         reg_in_n314, reg_in_n313, reg_in_n312, reg_in_n311, reg_in_n310,
         reg_in_n309, reg_in_n308, reg_in_n307, reg_in_n306, reg_in_n305,
         reg_in_n304, reg_in_n303, reg_in_n302, reg_in_n301, reg_in_n300,
         reg_in_n299, reg_in_n298, reg_in_n297, reg_in_n296, reg_in_n295,
         reg_in_n294, reg_in_n293, reg_in_n292, reg_in_n291, reg_in_n290,
         reg_in_n289, reg_in_n288, reg_in_n287, reg_in_n286, reg_in_n285,
         reg_in_n284, reg_in_n283, reg_in_n282, reg_in_n281, reg_in_n280,
         reg_in_n279, reg_in_n278, reg_in_n277, reg_in_n276, reg_in_n275,
         reg_in_n274, reg_in_n273, reg_in_n272, reg_in_n271, reg_in_n270,
         reg_in_n269, reg_in_n268, reg_in_n267, reg_in_n266, reg_in_n265,
         reg_in_n264, reg_in_n263, reg_in_n262, reg_in_n261, reg_in_n260,
         reg_in_n258, reg_in_n1, reg_in_pf0, reg_in_pf1, reg_in_pbv0,
         reg_in_pbv1, reg_out_n310, reg_out_n309, reg_out_n308, reg_out_n307,
         reg_out_n306, reg_out_n305, reg_out_n304, reg_out_n303, reg_out_n302,
         reg_out_n301, reg_out_n300, reg_out_n299, reg_out_n298, reg_out_n297,
         reg_out_n296, reg_out_n295, reg_out_n294, reg_out_n293, reg_out_n292,
         reg_out_n291, reg_out_n290, reg_out_n289, reg_out_n288, reg_out_n287,
         reg_out_n286, reg_out_n285, reg_out_n284, reg_out_n283, reg_out_n282,
         reg_out_n281, reg_out_n280, reg_out_n279, reg_out_n278, reg_out_n13,
         reg_out_n10, reg_out_n9, reg_out_n8, reg_out_n7, reg_out_n6,
         reg_out_n5, reg_out_n4, reg_out_n3, reg_out_n2, reg_out_n1,
         reg_out_n277, reg_out_n276, reg_out_n275, reg_out_n274, reg_out_n273,
         reg_out_n272, reg_out_n271, reg_out_n270, reg_out_n269, reg_out_n268,
         reg_out_n267, reg_out_n266, reg_out_n265, reg_out_n264, reg_out_n263,
         reg_out_n262, reg_out_n261, reg_out_n260, reg_out_n259, reg_out_n258,
         reg_out_n257, reg_out_n256, reg_out_n255, reg_out_n254, reg_out_n253,
         reg_out_n252, reg_out_n251, reg_out_n250, reg_out_n249, reg_out_n248,
         reg_out_n247, reg_out_n246, reg_out_n245, reg_out_n244, reg_out_n243,
         reg_out_n242, reg_out_n241, reg_out_n240, reg_out_n239, reg_out_n238,
         reg_out_n237, reg_out_n236, reg_out_n235, reg_out_n234, reg_out_n233,
         reg_out_n232, reg_out_n231, reg_out_n230, reg_out_n229, reg_out_n228,
         reg_out_n227, reg_out_n226, reg_out_n225, reg_out_n224, reg_out_n223,
         reg_out_n222, reg_out_n221, reg_out_n220, reg_out_n219, reg_out_n218,
         reg_out_n217, reg_out_n216, reg_out_n215, reg_out_n214, reg_out_n213,
         reg_out_n212, reg_out_n211, reg_out_n210, reg_out_n209, reg_out_n208,
         reg_out_n207, reg_out_n206, reg_out_n205, reg_out_n204, reg_out_n203,
         reg_out_n202, reg_out_n201, reg_out_n200, reg_out_n199, reg_out_n198,
         reg_out_n197, reg_out_n196, reg_out_n195, reg_out_n194, reg_out_n193,
         reg_out_n192, reg_out_n191, reg_out_n190, reg_out_n189, reg_out_n188,
         reg_out_n187, reg_out_n186, reg_out_n185, reg_out_n184, reg_out_n183,
         reg_out_n182, reg_out_n181, reg_out_n180, reg_out_n179, reg_out_n178,
         reg_out_n177, reg_out_n176, reg_out_n175, reg_out_n174, reg_out_n173,
         reg_out_n172, reg_out_n171, reg_out_n170, reg_out_n169, reg_out_n168,
         reg_out_n167, reg_out_n166, reg_out_n165, reg_out_n164, reg_out_n163,
         reg_out_n162, reg_out_n161, reg_out_n160, reg_out_n159, reg_out_n158,
         reg_out_n157, reg_out_n156, reg_out_n155, reg_out_n154, reg_out_n153,
         reg_out_n152, reg_out_n151, reg_out_n150, reg_out_n149, reg_out_n148,
         reg_out_n147, reg_out_n146, reg_out_n145, reg_out_n144, reg_out_n143,
         reg_out_n142, reg_out_n141, reg_out_n140, reg_out_n139, reg_out_n138,
         reg_out_n137, reg_out_n136, reg_out_n135, reg_out_n134, reg_out_n133,
         reg_out_n132, reg_out_n131, reg_out_n130, reg_out_n129, reg_out_n128,
         reg_out_n127, reg_out_n126, reg_out_n125, reg_out_n124, reg_out_n123,
         reg_out_n122, reg_out_n121, reg_out_n120, reg_out_n119, reg_out_n118,
         reg_out_n117, reg_out_n116, reg_out_n115, reg_out_n114, reg_out_n113,
         reg_out_n112, reg_out_n111, reg_out_n110, reg_out_n109, reg_out_n108,
         reg_out_n107, reg_out_n106, reg_out_n105, reg_out_n104, reg_out_n103,
         reg_out_n102, reg_out_n101, reg_out_n100, reg_out_n99, reg_out_n98,
         reg_out_n97, reg_out_n96, reg_out_n95, reg_out_n94, reg_out_n93,
         reg_out_n92, reg_out_n91, reg_out_n90, reg_out_n89, reg_out_n88,
         reg_out_n87, reg_out_n86, reg_out_n85, reg_out_n84, reg_out_n83,
         reg_out_n82, reg_out_n81, reg_out_n80, reg_out_n79, reg_out_n78,
         reg_out_n77, reg_out_n76, reg_out_n75, reg_out_n74, reg_out_n73,
         reg_out_n72, reg_out_n71, reg_out_n70, reg_out_n69, reg_out_n68,
         reg_out_n67, reg_out_n66, reg_out_n65, reg_out_n64, reg_out_n63,
         reg_out_n62, reg_out_n61, reg_out_n60, reg_out_n59, reg_out_n58,
         reg_out_n57, reg_out_n56, reg_out_n55, reg_out_n54, reg_out_n53,
         reg_out_n52, reg_out_n51, reg_out_n50, reg_out_n49, reg_out_n48,
         reg_out_n47, reg_out_n46, reg_out_n45, reg_out_n44, reg_out_n43,
         reg_out_n42, reg_out_n41, reg_out_n40, reg_out_n39, reg_out_n38,
         reg_out_n37, reg_out_n36, reg_out_n35, reg_out_n34, reg_out_n33,
         reg_out_n32, reg_out_n31, reg_out_n30, reg_out_n29, reg_out_n28,
         reg_out_n27, reg_out_n26, reg_out_n25, reg_out_n24, reg_out_n23,
         reg_out_n22, reg_out_n21, reg_out_n20, reg_out_n19, reg_out_n18,
         reg_out_n17, reg_out_n16, reg_out_n15, reg_out_n14, reg_out_n12,
         reg_out_n11, reg_out_rdy1, reg_out_rdy2, reg_out_rdy0;
  wire   [255:0] Din;
  wire   [127:0] Dout;
  wire   [6:0] control_gray_dout;
  wire   [6:0] control_bin_add;
  wire   [6:0] control_bin_dout;
  wire   [6:2] control_add_15_carry;
  wire   [1:0] aes_core_aes_core_ctrl_reg;
  wire   [31:0] aes_core_keymem_sboxw;
  wire   [31:0] aes_core_new_sboxw;
  wire   [31:0] aes_core_enc_sboxw;
  wire   [127:0] aes_core_round_key;
  wire   [3:0] aes_core_enc_round_nr;
  wire   [1:0] aes_core_enc_block_enc_ctrl_reg;
  wire   [1:0] aes_core_enc_block_sword_ctr_reg;
  wire   [127:32] aes_core_keymem_prev_key1_reg;
  wire   [1407:0] aes_core_keymem_key_mem;
  wire   [3:0] aes_core_keymem_round_ctr_reg;
  wire   [1:0] aes_core_keymem_key_mem_ctrl_reg;
  wire   [7:0] aes_core_keymem_rcon_reg;
  wire   [255:0] reg_in_plain_text;
  wire   [127:0] reg_out_cipher_sample;
  CLKINVX4 U1 ( .A(reset_p), .Y(reset_n) );
  XNOR2X1 control_U30 ( .A(control_gray_dout[0]), .B(control_gray_dout[3]), 
        .Y(control_n5) );
  NOR3X1 control_U29 ( .A(control_gray_dout[1]), .B(control_gray_dout[6]), .C(
        control_gray_dout[5]), .Y(control_n6) );
  NAND4X1 control_U28 ( .A(control_gray_dout[4]), .B(control_gray_dout[2]), 
        .C(control_n5), .D(control_n6), .Y(control_n4) );
  OAI2BB2X1 control_U27 ( .B0(control_n3), .B1(control_n4), .A0N(next), .A1N(
        control_n4), .Y(control_n19) );
  INVX1 control_U26 ( .A(control_gray_dout[3]), .Y(control_n2) );
  NAND3BX1 control_U25 ( .AN(control_gray_dout[2]), .B(control_n2), .C(
        control_n8), .Y(control_n9) );
  OAI2BB2X1 control_U24 ( .B0(control_n1), .B1(control_n9), .A0N(trig), .A1N(
        control_n9), .Y(control_n21) );
  NAND3X1 control_U23 ( .A(control_gray_dout[2]), .B(control_gray_dout[3]), 
        .C(control_n8), .Y(control_n7) );
  OAI2BB2X1 control_U22 ( .B0(control_n3), .B1(control_n7), .A0N(init), .A1N(
        control_n7), .Y(control_n20) );
  INVX1 control_U21 ( .A(control_gray_dout[0]), .Y(control_n1) );
  NAND3X1 control_U20 ( .A(control_gray_dout[0]), .B(control_gray_dout[3]), 
        .C(control_gray_dout[2]), .Y(control_n3) );
  XNOR2X1 control_U19 ( .A(control_gray_dout[1]), .B(control_n1), .Y(
        control_n10) );
  NOR4BX1 control_U18 ( .AN(control_n10), .B(control_gray_dout[4]), .C(
        control_gray_dout[5]), .D(control_gray_dout[6]), .Y(control_n8) );
  NOR2BX1 control_U17 ( .AN(control_gray_dout[4]), .B(control_n3), .Y(
        control_n18) );
  AND4X2 control_U16 ( .A(control_gray_dout[6]), .B(control_gray_dout[5]), .C(
        control_n18), .D(control_gray_dout[1]), .Y(control_n11) );
  XNOR2X1 control_U15 ( .A(control_bin_add[1]), .B(control_bin_add[0]), .Y(
        control_n17) );
  NOR2X1 control_U14 ( .A(control_n11), .B(control_n17), .Y(control_N100) );
  XNOR2X1 control_U13 ( .A(control_bin_add[1]), .B(control_bin_add[2]), .Y(
        control_n16) );
  NOR2X1 control_U12 ( .A(control_n11), .B(control_n16), .Y(control_N110) );
  XNOR2X1 control_U11 ( .A(control_bin_add[2]), .B(control_bin_add[3]), .Y(
        control_n15) );
  NOR2X1 control_U10 ( .A(control_n11), .B(control_n15), .Y(control_N120) );
  XNOR2X1 control_U9 ( .A(control_bin_add[3]), .B(control_bin_add[4]), .Y(
        control_n14) );
  NOR2X1 control_U8 ( .A(control_n11), .B(control_n14), .Y(control_N130) );
  NOR2BX1 control_U7 ( .AN(control_bin_add[6]), .B(control_n11), .Y(
        control_N160) );
  XNOR2X1 control_U6 ( .A(control_bin_add[4]), .B(control_bin_add[5]), .Y(
        control_n13) );
  NOR2X1 control_U5 ( .A(control_n11), .B(control_n13), .Y(control_N140) );
  XNOR2X1 control_U4 ( .A(control_bin_add[5]), .B(control_bin_add[6]), .Y(
        control_n12) );
  NOR2X1 control_U3 ( .A(control_n11), .B(control_n12), .Y(control_N150) );
  DFFRHQX1 control_trig_reg ( .D(control_n21), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(trig) );
  DFFRHQX1 control_init_reg ( .D(control_n20), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(init) );
  DFFRHQX1 control_next_reg ( .D(control_n19), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(next) );
  DFFRHQX1 control_gray_dout_reg_3_ ( .D(control_N130), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[3]) );
  DFFRHQX1 control_gray_dout_reg_6_ ( .D(control_N160), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[6]) );
  DFFRHQX1 control_gray_dout_reg_4_ ( .D(control_N140), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[4]) );
  DFFRHQX1 control_gray_dout_reg_5_ ( .D(control_N150), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[5]) );
  DFFRHQX1 control_gray_dout_reg_2_ ( .D(control_N120), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[2]) );
  DFFRHQX1 control_gray_dout_reg_1_ ( .D(control_N110), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[1]) );
  DFFRHQX1 control_gray_dout_reg_0_ ( .D(control_N100), .CK(clk_48Mhz), .RN(
        reset_n), .Q(control_gray_dout[0]) );
  BUFX3 control_gtb_U7 ( .A(control_gray_dout[6]), .Y(control_bin_dout[6]) );
  XOR2X1 control_gtb_U6 ( .A(control_gray_dout[0]), .B(control_bin_dout[1]), 
        .Y(control_bin_dout[0]) );
  XOR2X1 control_gtb_U5 ( .A(control_bin_dout[5]), .B(control_gray_dout[4]), 
        .Y(control_bin_dout[4]) );
  XOR2X1 control_gtb_U4 ( .A(control_bin_dout[3]), .B(control_gray_dout[2]), 
        .Y(control_bin_dout[2]) );
  XOR2X1 control_gtb_U3 ( .A(control_bin_dout[4]), .B(control_gray_dout[3]), 
        .Y(control_bin_dout[3]) );
  XOR2X1 control_gtb_U2 ( .A(control_gray_dout[5]), .B(control_gray_dout[6]), 
        .Y(control_bin_dout[5]) );
  XOR2X1 control_gtb_U1 ( .A(control_bin_dout[2]), .B(control_gray_dout[1]), 
        .Y(control_bin_dout[1]) );
  INVX1 control_add_15_U2 ( .A(control_bin_dout[0]), .Y(control_bin_add[0]) );
  XOR2X1 control_add_15_U1 ( .A(control_add_15_carry[6]), .B(
        control_bin_dout[6]), .Y(control_bin_add[6]) );
  CMPR22X1 control_add_15_U1_1_1 ( .A(control_bin_dout[1]), .B(
        control_bin_dout[0]), .CO(control_add_15_carry[2]), .S(
        control_bin_add[1]) );
  CMPR22X1 control_add_15_U1_1_2 ( .A(control_bin_dout[2]), .B(
        control_add_15_carry[2]), .CO(control_add_15_carry[3]), .S(
        control_bin_add[2]) );
  CMPR22X1 control_add_15_U1_1_3 ( .A(control_bin_dout[3]), .B(
        control_add_15_carry[3]), .CO(control_add_15_carry[4]), .S(
        control_bin_add[3]) );
  CMPR22X1 control_add_15_U1_1_4 ( .A(control_bin_dout[4]), .B(
        control_add_15_carry[4]), .CO(control_add_15_carry[5]), .S(
        control_bin_add[4]) );
  CMPR22X1 control_add_15_U1_1_5 ( .A(control_bin_dout[5]), .B(
        control_add_15_carry[5]), .CO(control_add_15_carry[6]), .S(
        control_bin_add[5]) );
  OAI2BB1X1 aes_core_U95 ( .A0N(ready), .A1N(aes_core_n38), .B0(aes_core_n39), 
        .Y(aes_core_n75) );
  INVX1 aes_core_U94 ( .A(aes_core_aes_core_ctrl_reg[1]), .Y(aes_core_n92) );
  AOI2BB1X1 aes_core_U93 ( .A0N(init), .A1N(next), .B0(aes_core_n40), .Y(
        aes_core_n41) );
  NOR2BX1 aes_core_U92 ( .AN(aes_core_n39), .B(aes_core_n41), .Y(aes_core_n38)
         );
  OAI32X1 aes_core_U91 ( .A0(aes_core_n40), .A1(init), .A2(aes_core_n38), .B0(
        aes_core_n92), .B1(aes_core_n90), .Y(aes_core_n76) );
  AOI33X1 aes_core_U90 ( .A0(aes_core_aes_core_ctrl_reg[1]), .A1(aes_core_n91), 
        .A2(aes_core_enc_ready), .B0(aes_core_aes_core_ctrl_reg[0]), .B1(
        aes_core_n92), .B2(aes_core_key_ready), .Y(aes_core_n39) );
  AOI22X1 aes_core_U89 ( .A0(aes_core_enc_sboxw[31]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[31]), .B1(aes_core_n80), .Y(aes_core_n50) );
  INVX1 aes_core_U88 ( .A(aes_core_n50), .Y(aes_core_n33) );
  AOI22X1 aes_core_U87 ( .A0(aes_core_enc_sboxw[23]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[23]), .B1(aes_core_n80), .Y(aes_core_n59) );
  INVX1 aes_core_U86 ( .A(aes_core_n59), .Y(aes_core_n25) );
  AOI22X1 aes_core_U85 ( .A0(aes_core_enc_sboxw[22]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[22]), .B1(aes_core_n81), .Y(aes_core_n60) );
  INVX1 aes_core_U84 ( .A(aes_core_n60), .Y(aes_core_n24) );
  AOI22X1 aes_core_U83 ( .A0(aes_core_enc_sboxw[15]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[15]), .B1(aes_core_n84), .Y(aes_core_n68) );
  INVX1 aes_core_U82 ( .A(aes_core_n68), .Y(aes_core_n17) );
  AOI22X1 aes_core_U81 ( .A0(aes_core_enc_sboxw[7]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[7]), .B1(aes_core_n34), .Y(aes_core_n45) );
  INVX1 aes_core_U80 ( .A(aes_core_n45), .Y(aes_core_n9) );
  AOI22X1 aes_core_U79 ( .A0(aes_core_enc_sboxw[14]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[14]), .B1(aes_core_n83), .Y(aes_core_n69) );
  INVX1 aes_core_U78 ( .A(aes_core_n69), .Y(aes_core_n16) );
  AOI22X1 aes_core_U77 ( .A0(aes_core_enc_sboxw[6]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[6]), .B1(aes_core_n83), .Y(aes_core_n46) );
  INVX1 aes_core_U76 ( .A(aes_core_n46), .Y(aes_core_n8) );
  AOI22X1 aes_core_U75 ( .A0(aes_core_enc_sboxw[30]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[30]), .B1(aes_core_n81), .Y(aes_core_n51) );
  INVX1 aes_core_U74 ( .A(aes_core_n51), .Y(aes_core_n32) );
  INVX1 aes_core_U73 ( .A(aes_core_aes_core_ctrl_reg[0]), .Y(aes_core_n91) );
  AOI22X1 aes_core_U72 ( .A0(aes_core_enc_sboxw[29]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[29]), .B1(aes_core_n82), .Y(aes_core_n53) );
  INVX1 aes_core_U71 ( .A(aes_core_n53), .Y(aes_core_n31) );
  AOI22X1 aes_core_U70 ( .A0(aes_core_enc_sboxw[26]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[26]), .B1(aes_core_n82), .Y(aes_core_n56) );
  INVX1 aes_core_U69 ( .A(aes_core_n56), .Y(aes_core_n28) );
  AOI22X1 aes_core_U68 ( .A0(aes_core_enc_sboxw[12]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[12]), .B1(aes_core_n85), .Y(aes_core_n71) );
  AOI22X1 aes_core_U67 ( .A0(aes_core_enc_sboxw[28]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[28]), .B1(aes_core_n84), .Y(aes_core_n54) );
  AOI22X1 aes_core_U66 ( .A0(aes_core_enc_sboxw[5]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[5]), .B1(aes_core_n80), .Y(aes_core_n47) );
  INVX1 aes_core_U65 ( .A(aes_core_n47), .Y(aes_core_n7) );
  AOI22X1 aes_core_U64 ( .A0(aes_core_enc_sboxw[21]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[21]), .B1(aes_core_n82), .Y(aes_core_n61) );
  INVX1 aes_core_U63 ( .A(aes_core_n61), .Y(aes_core_n23) );
  AOI22X1 aes_core_U62 ( .A0(aes_core_enc_sboxw[0]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[0]), .B1(aes_core_n85), .Y(aes_core_n74) );
  INVX1 aes_core_U61 ( .A(aes_core_n74), .Y(aes_core_n2) );
  AOI22X1 aes_core_U60 ( .A0(aes_core_enc_sboxw[1]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[1]), .B1(aes_core_n83), .Y(aes_core_n63) );
  INVX1 aes_core_U59 ( .A(aes_core_n63), .Y(aes_core_n3) );
  AOI22X1 aes_core_U58 ( .A0(aes_core_enc_sboxw[16]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[16]), .B1(aes_core_n84), .Y(aes_core_n67) );
  INVX1 aes_core_U57 ( .A(aes_core_n67), .Y(aes_core_n18) );
  AOI22X1 aes_core_U56 ( .A0(aes_core_enc_sboxw[17]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[17]), .B1(aes_core_n83), .Y(aes_core_n66) );
  INVX1 aes_core_U55 ( .A(aes_core_n66), .Y(aes_core_n19) );
  AOI22X1 aes_core_U54 ( .A0(aes_core_enc_sboxw[24]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[24]), .B1(aes_core_n84), .Y(aes_core_n58) );
  INVX1 aes_core_U53 ( .A(aes_core_n58), .Y(aes_core_n26) );
  AOI22X1 aes_core_U52 ( .A0(aes_core_enc_sboxw[25]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[25]), .B1(aes_core_n82), .Y(aes_core_n57) );
  INVX1 aes_core_U51 ( .A(aes_core_n57), .Y(aes_core_n27) );
  AOI22X1 aes_core_U50 ( .A0(aes_core_enc_sboxw[10]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[10]), .B1(aes_core_n85), .Y(aes_core_n73) );
  AOI22X1 aes_core_U49 ( .A0(aes_core_enc_sboxw[11]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[11]), .B1(aes_core_n83), .Y(aes_core_n72) );
  INVX1 aes_core_U48 ( .A(aes_core_n72), .Y(aes_core_n13) );
  AOI22X1 aes_core_U47 ( .A0(aes_core_enc_sboxw[27]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[27]), .B1(aes_core_n82), .Y(aes_core_n55) );
  INVX1 aes_core_U46 ( .A(aes_core_n55), .Y(aes_core_n29) );
  AOI22X1 aes_core_U45 ( .A0(aes_core_enc_sboxw[19]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[19]), .B1(aes_core_n83), .Y(aes_core_n64) );
  INVX1 aes_core_U44 ( .A(aes_core_n64), .Y(aes_core_n21) );
  INVX1 aes_core_U43 ( .A(aes_core_n38), .Y(aes_core_n90) );
  OAI22X1 aes_core_U42 ( .A0(aes_core_n91), .A1(aes_core_n90), .B0(
        aes_core_n40), .B1(aes_core_n93), .Y(aes_core_n77) );
  NAND2X1 aes_core_U41 ( .A(aes_core_n91), .B(aes_core_n92), .Y(aes_core_n40)
         );
  INVX1 aes_core_U40 ( .A(aes_core_n43), .Y(aes_core_n35) );
  INVX1 aes_core_U39 ( .A(aes_core_n43), .Y(aes_core_n36) );
  INVX1 aes_core_U38 ( .A(aes_core_n36), .Y(aes_core_n1) );
  INVX1 aes_core_U37 ( .A(aes_core_n85), .Y(aes_core_n89) );
  INVX1 aes_core_U36 ( .A(aes_core_n34), .Y(aes_core_n88) );
  INVX1 aes_core_U35 ( .A(aes_core_n87), .Y(aes_core_n85) );
  INVX1 aes_core_U34 ( .A(aes_core_n89), .Y(aes_core_n84) );
  INVX1 aes_core_U33 ( .A(aes_core_n87), .Y(aes_core_n86) );
  INVX1 aes_core_U32 ( .A(aes_core_n89), .Y(aes_core_n81) );
  INVX1 aes_core_U31 ( .A(aes_core_n89), .Y(aes_core_n80) );
  INVX1 aes_core_U30 ( .A(aes_core_n88), .Y(aes_core_n82) );
  AOI22X2 aes_core_U29 ( .A0(aes_core_enc_sboxw[2]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[2]), .B1(aes_core_n81), .Y(aes_core_n52) );
  AOI22X2 aes_core_U28 ( .A0(aes_core_enc_sboxw[20]), .A1(aes_core_n78), .B0(
        aes_core_keymem_sboxw[20]), .B1(aes_core_n82), .Y(aes_core_n62) );
  AOI22X4 aes_core_U27 ( .A0(aes_core_enc_sboxw[9]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[9]), .B1(aes_core_n82), .Y(aes_core_n42) );
  AOI22X4 aes_core_U26 ( .A0(aes_core_enc_sboxw[3]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[3]), .B1(aes_core_n81), .Y(aes_core_n49) );
  AOI22X1 aes_core_U25 ( .A0(aes_core_enc_sboxw[18]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[18]), .B1(aes_core_n83), .Y(aes_core_n65) );
  INVX1 aes_core_U24 ( .A(aes_core_n65), .Y(aes_core_n20) );
  AOI22X1 aes_core_U23 ( .A0(aes_core_enc_sboxw[13]), .A1(aes_core_n37), .B0(
        aes_core_keymem_sboxw[13]), .B1(aes_core_n82), .Y(aes_core_n70) );
  INVX1 aes_core_U22 ( .A(aes_core_n70), .Y(aes_core_n15) );
  CLKINVX8 aes_core_U21 ( .A(aes_core_n49), .Y(aes_core_n5) );
  CLKINVX8 aes_core_U20 ( .A(aes_core_n48), .Y(aes_core_n6) );
  CLKINVX8 aes_core_U19 ( .A(aes_core_n62), .Y(aes_core_n22) );
  CLKINVX8 aes_core_U18 ( .A(aes_core_n52), .Y(aes_core_n4) );
  INVX1 aes_core_U17 ( .A(aes_core_n88), .Y(aes_core_n83) );
  INVX4 aes_core_U16 ( .A(aes_core_n1), .Y(aes_core_n87) );
  INVX1 aes_core_U15 ( .A(aes_core_n73), .Y(aes_core_n12) );
  INVX8 aes_core_U14 ( .A(aes_core_n42), .Y(aes_core_n11) );
  INVX1 aes_core_U13 ( .A(aes_core_n35), .Y(aes_core_n34) );
  INVX1 aes_core_U12 ( .A(aes_core_n86), .Y(aes_core_n79) );
  INVX1 aes_core_U11 ( .A(aes_core_n86), .Y(aes_core_n78) );
  AOI22X1 aes_core_U10 ( .A0(aes_core_enc_sboxw[8]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[8]), .B1(aes_core_n82), .Y(aes_core_n44) );
  INVX1 aes_core_U9 ( .A(aes_core_n44), .Y(aes_core_n10) );
  CLKINVX4 aes_core_U8 ( .A(aes_core_n71), .Y(aes_core_n14) );
  CLKINVX3 aes_core_U7 ( .A(aes_core_n86), .Y(aes_core_n37) );
  INVX1 aes_core_U6 ( .A(init), .Y(aes_core_n93) );
  AOI21X1 aes_core_U5 ( .A0(aes_core_n93), .A1(aes_core_n91), .B0(
        aes_core_aes_core_ctrl_reg[1]), .Y(aes_core_n43) );
  CLKINVX3 aes_core_U4 ( .A(aes_core_n54), .Y(aes_core_n30) );
  AOI22X1 aes_core_U3 ( .A0(aes_core_enc_sboxw[4]), .A1(aes_core_n79), .B0(
        aes_core_keymem_sboxw[4]), .B1(aes_core_n80), .Y(aes_core_n48) );
  DFFRHQX1 aes_core_aes_core_ctrl_reg_reg_0_ ( .D(aes_core_n77), .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_aes_core_ctrl_reg[0]) );
  DFFRHQX1 aes_core_aes_core_ctrl_reg_reg_1_ ( .D(aes_core_n76), .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_aes_core_ctrl_reg[1]) );
  DFFSX1 aes_core_ready_reg_reg ( .D(aes_core_n75), .CK(clk_48Mhz), .SN(
        reset_n), .Q(ready), .QN() );
  DFFRX1 aes_core_enc_block_block_w1_reg_reg_0_ ( .D(aes_core_enc_block_n1273), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[64]), .QN(
        aes_core_enc_block_n1362) );
  OAI22X1 aes_core_enc_block_U1492 ( .A0(aes_core_enc_block_n182), .A1(
        aes_core_enc_block_n1205), .B0(aes_core_enc_round_nr[0]), .B1(
        aes_core_enc_block_n1203), .Y(aes_core_enc_block_n1342) );
  INVX1 aes_core_enc_block_U1491 ( .A(Dout[27]), .Y(aes_core_enc_block_n1451)
         );
  NAND3X1 aes_core_enc_block_U1490 ( .A(aes_core_enc_block_n180), .B(
        aes_core_enc_block_n181), .C(next), .Y(aes_core_enc_block_n1196) );
  INVX1 aes_core_enc_block_U1489 ( .A(Dout[7]), .Y(aes_core_enc_block_n1384)
         );
  INVX1 aes_core_enc_block_U1488 ( .A(Dout[12]), .Y(aes_core_enc_block_n1351)
         );
  INVX1 aes_core_enc_block_U1487 ( .A(Dout[26]), .Y(aes_core_enc_block_n1447)
         );
  INVX1 aes_core_enc_block_U1486 ( .A(Dout[40]), .Y(aes_core_enc_block_n1423)
         );
  INVX1 aes_core_enc_block_U1485 ( .A(Dout[56]), .Y(aes_core_enc_block_n1395)
         );
  INVX1 aes_core_enc_block_U1484 ( .A(Dout[24]), .Y(aes_core_enc_block_n1425)
         );
  INVX1 aes_core_enc_block_U1483 ( .A(Dout[14]), .Y(aes_core_enc_block_n1381)
         );
  INVX1 aes_core_enc_block_U1482 ( .A(Dout[13]), .Y(aes_core_enc_block_n1369)
         );
  INVX1 aes_core_enc_block_U1481 ( .A(aes_core_enc_round_nr[0]), .Y(
        aes_core_enc_block_n182) );
  INVX1 aes_core_enc_block_U1480 ( .A(Dout[29]), .Y(aes_core_enc_block_n1379)
         );
  INVX1 aes_core_enc_block_U1479 ( .A(Dout[30]), .Y(aes_core_enc_block_n1380)
         );
  OAI2BB1X1 aes_core_enc_block_U1478 ( .A0N(aes_core_enc_ready), .A1N(
        aes_core_enc_block_n1196), .B0(aes_core_enc_block_n81), .Y(
        aes_core_enc_block_n1339) );
  AOI32X1 aes_core_enc_block_U1477 ( .A0(aes_core_enc_round_nr[1]), .A1(
        aes_core_enc_block_n185), .A2(aes_core_enc_block_n1200), .B0(
        aes_core_enc_block_n1201), .B1(aes_core_enc_round_nr[2]), .Y(
        aes_core_enc_block_n1202) );
  INVX1 aes_core_enc_block_U1476 ( .A(aes_core_enc_block_n1202), .Y(
        aes_core_enc_block_n175) );
  AOI21X1 aes_core_enc_block_U1475 ( .A0(aes_core_enc_block_n177), .A1(
        aes_core_enc_block_n185), .B0(aes_core_enc_block_n1201), .Y(
        aes_core_enc_block_n1198) );
  NAND4X1 aes_core_enc_block_U1474 ( .A(aes_core_enc_round_nr[2]), .B(
        aes_core_enc_round_nr[1]), .C(aes_core_enc_block_n1200), .D(
        aes_core_enc_block_n186), .Y(aes_core_enc_block_n1199) );
  OAI21X1 aes_core_enc_block_U1473 ( .A0(aes_core_enc_block_n1198), .A1(
        aes_core_enc_block_n186), .B0(aes_core_enc_block_n1199), .Y(
        aes_core_enc_block_n1340) );
  XNOR2X1 aes_core_enc_block_U1472 ( .A(aes_core_enc_block_n1364), .B(Dout[66]), .Y(aes_core_enc_block_n759) );
  XNOR2X1 aes_core_enc_block_U1471 ( .A(aes_core_enc_block_n1412), .B(Dout[94]), .Y(aes_core_enc_block_n475) );
  XNOR2X1 aes_core_enc_block_U1470 ( .A(aes_core_enc_block_n1454), .B(Dout[74]), .Y(aes_core_enc_block_n998) );
  XNOR2X1 aes_core_enc_block_U1469 ( .A(aes_core_enc_block_n1449), .B(Dout[83]), .Y(aes_core_enc_block_n267) );
  XNOR2X1 aes_core_enc_block_U1468 ( .A(aes_core_enc_block_n1458), .B(Dout[98]), .Y(aes_core_enc_block_n518) );
  XNOR2X1 aes_core_enc_block_U1467 ( .A(aes_core_enc_block_n1356), .B(Dout[6]), 
        .Y(aes_core_enc_block_n251) );
  XNOR2X1 aes_core_enc_block_U1466 ( .A(aes_core_enc_block_n1375), .B(Dout[99]), .Y(aes_core_enc_block_n509) );
  XNOR2X1 aes_core_enc_block_U1465 ( .A(aes_core_enc_block_n190), .B(Dout[67]), 
        .Y(aes_core_enc_block_n750) );
  XNOR2X1 aes_core_enc_block_U1464 ( .A(aes_core_enc_block_n191), .B(Dout[75]), 
        .Y(aes_core_enc_block_n989) );
  XNOR2X1 aes_core_enc_block_U1463 ( .A(aes_core_enc_block_n1421), .B(Dout[80]), .Y(aes_core_enc_block_n295) );
  XNOR2X1 aes_core_enc_block_U1462 ( .A(aes_core_enc_block_n1457), .B(Dout[42]), .Y(aes_core_enc_block_n286) );
  XNOR2X1 aes_core_enc_block_U1461 ( .A(aes_core_enc_block_n1409), .B(Dout[86]), .Y(aes_core_enc_block_n243) );
  XNOR2X1 aes_core_enc_block_U1460 ( .A(aes_core_enc_block_n1365), .B(Dout[91]), .Y(aes_core_enc_block_n499) );
  XNOR2X1 aes_core_enc_block_U1459 ( .A(aes_core_enc_block_n1411), .B(Dout[62]), .Y(aes_core_enc_block_n716) );
  XNOR2X1 aes_core_enc_block_U1458 ( .A(aes_core_enc_block_n1410), .B(Dout[30]), .Y(aes_core_enc_block_n955) );
  XNOR2X1 aes_core_enc_block_U1457 ( .A(aes_core_enc_block_n232), .B(Dout[78]), 
        .Y(aes_core_enc_block_n963) );
  XNOR2X1 aes_core_enc_block_U1456 ( .A(aes_core_enc_block_n1455), .B(Dout[43]), .Y(aes_core_enc_block_n277) );
  XNOR2X1 aes_core_enc_block_U1455 ( .A(aes_core_enc_block_n196), .B(Dout[70]), 
        .Y(aes_core_enc_block_n724) );
  XNOR2X1 aes_core_enc_block_U1454 ( .A(aes_core_enc_block_n1427), .B(Dout[88]), .Y(aes_core_enc_block_n527) );
  XNOR2X1 aes_core_enc_block_U1453 ( .A(aes_core_enc_block_n1357), .B(Dout[14]), .Y(aes_core_enc_block_n483) );
  XNOR2X1 aes_core_enc_block_U1452 ( .A(aes_core_enc_block_n1400), .B(Dout[59]), .Y(aes_core_enc_block_n740) );
  XNOR2X1 aes_core_enc_block_U1451 ( .A(aes_core_enc_block_n1424), .B(Dout[24]), .Y(aes_core_enc_block_n1007) );
  XNOR2X1 aes_core_enc_block_U1450 ( .A(aes_core_enc_block_n1426), .B(Dout[56]), .Y(aes_core_enc_block_n768) );
  XNOR2X1 aes_core_enc_block_U1449 ( .A(aes_core_enc_block_n1450), .B(Dout[27]), .Y(aes_core_enc_block_n979) );
  OAI21X1 aes_core_enc_block_U1448 ( .A0(aes_core_enc_block_n1203), .A1(
        aes_core_enc_round_nr[1]), .B0(aes_core_enc_block_n1204), .Y(
        aes_core_enc_block_n1201) );
  XNOR2X1 aes_core_enc_block_U1447 ( .A(aes_core_enc_block_n1406), .B(Dout[93]), .Y(aes_core_enc_block_n484) );
  XNOR2X1 aes_core_enc_block_U1446 ( .A(aes_core_enc_block_n1401), .B(Dout[92]), .Y(aes_core_enc_block_n492) );
  XNOR2X1 aes_core_enc_block_U1445 ( .A(aes_core_enc_block_n1353), .B(Dout[5]), 
        .Y(aes_core_enc_block_n259) );
  XNOR2X1 aes_core_enc_block_U1444 ( .A(aes_core_enc_block_n1445), .B(Dout[82]), .Y(aes_core_enc_block_n278) );
  XNOR2X1 aes_core_enc_block_U1443 ( .A(aes_core_enc_block_n1387), .B(Dout[84]), .Y(aes_core_enc_block_n260) );
  XNOR2X1 aes_core_enc_block_U1442 ( .A(aes_core_enc_block_n1434), .B(Dout[81]), .Y(aes_core_enc_block_n287) );
  XNOR2X1 aes_core_enc_block_U1441 ( .A(aes_core_enc_block_n194), .B(Dout[77]), 
        .Y(aes_core_enc_block_n971) );
  XNOR2X1 aes_core_enc_block_U1440 ( .A(aes_core_enc_block_n1436), .B(Dout[65]), .Y(aes_core_enc_block_n767) );
  XNOR2X1 aes_core_enc_block_U1439 ( .A(aes_core_enc_block_n1349), .B(Dout[68]), .Y(aes_core_enc_block_n742) );
  XNOR2X1 aes_core_enc_block_U1438 ( .A(aes_core_enc_block_n1396), .B(Dout[72]), .Y(aes_core_enc_block_n1015) );
  XNOR2X1 aes_core_enc_block_U1437 ( .A(aes_core_enc_block_n1422), .B(Dout[64]), .Y(aes_core_enc_block_n776) );
  XNOR2X1 aes_core_enc_block_U1436 ( .A(aes_core_enc_block_n1377), .B(Dout[4]), 
        .Y(aes_core_enc_block_n269) );
  XNOR2X1 aes_core_enc_block_U1435 ( .A(aes_core_enc_block_n1397), .B(Dout[41]), .Y(aes_core_enc_block_n294) );
  XNOR2X1 aes_core_enc_block_U1434 ( .A(aes_core_enc_block_n1350), .B(Dout[76]), .Y(aes_core_enc_block_n981) );
  XNOR2X1 aes_core_enc_block_U1433 ( .A(aes_core_enc_block_n1456), .B(Dout[73]), .Y(aes_core_enc_block_n1006) );
  XNOR2X1 aes_core_enc_block_U1432 ( .A(aes_core_enc_block_n1408), .B(Dout[85]), .Y(aes_core_enc_block_n252) );
  XNOR2X1 aes_core_enc_block_U1431 ( .A(aes_core_enc_block_n1442), .B(Dout[90]), .Y(aes_core_enc_block_n510) );
  XNOR2X1 aes_core_enc_block_U1430 ( .A(aes_core_enc_block_n1431), .B(Dout[89]), .Y(aes_core_enc_block_n519) );
  XNOR2X1 aes_core_enc_block_U1429 ( .A(aes_core_enc_block_n1405), .B(Dout[61]), .Y(aes_core_enc_block_n725) );
  XNOR2X1 aes_core_enc_block_U1428 ( .A(aes_core_enc_block_n1378), .B(Dout[29]), .Y(aes_core_enc_block_n964) );
  XNOR2X1 aes_core_enc_block_U1427 ( .A(aes_core_enc_block_n1390), .B(Dout[60]), .Y(aes_core_enc_block_n733) );
  XNOR2X1 aes_core_enc_block_U1426 ( .A(aes_core_enc_block_n1439), .B(Dout[57]), .Y(aes_core_enc_block_n760) );
  XNOR2X1 aes_core_enc_block_U1425 ( .A(aes_core_enc_block_n193), .B(Dout[69]), 
        .Y(aes_core_enc_block_n732) );
  XNOR2X1 aes_core_enc_block_U1424 ( .A(aes_core_enc_block_n947), .B(Dout[40]), 
        .Y(aes_core_enc_block_n303) );
  XNOR2X1 aes_core_enc_block_U1423 ( .A(aes_core_enc_block_n1428), .B(Dout[96]), .Y(aes_core_enc_block_n535) );
  XNOR2X1 aes_core_enc_block_U1422 ( .A(aes_core_enc_block_n1354), .B(Dout[13]), .Y(aes_core_enc_block_n491) );
  XNOR2X1 aes_core_enc_block_U1421 ( .A(aes_core_enc_block_n1448), .B(Dout[58]), .Y(aes_core_enc_block_n751) );
  XNOR2X1 aes_core_enc_block_U1420 ( .A(aes_core_enc_block_n1388), .B(Dout[28]), .Y(aes_core_enc_block_n972) );
  XNOR2X1 aes_core_enc_block_U1419 ( .A(aes_core_enc_block_n1435), .B(Dout[25]), .Y(aes_core_enc_block_n999) );
  XNOR2X1 aes_core_enc_block_U1418 ( .A(aes_core_enc_block_n1446), .B(Dout[26]), .Y(aes_core_enc_block_n990) );
  XNOR2X1 aes_core_enc_block_U1417 ( .A(aes_core_enc_block_n1367), .B(Dout[12]), .Y(aes_core_enc_block_n501) );
  XNOR2X1 aes_core_enc_block_U1416 ( .A(aes_core_enc_block_n1207), .B(Dout[9]), 
        .Y(aes_core_enc_block_n526) );
  INVX1 aes_core_enc_block_U1415 ( .A(Dout[11]), .Y(aes_core_enc_block_n1375)
         );
  INVX1 aes_core_enc_block_U1414 ( .A(Dout[51]), .Y(aes_core_enc_block_n1365)
         );
  INVX1 aes_core_enc_block_U1413 ( .A(Dout[48]), .Y(aes_core_enc_block_n1427)
         );
  INVX1 aes_core_enc_block_U1412 ( .A(Dout[50]), .Y(aes_core_enc_block_n1442)
         );
  INVX1 aes_core_enc_block_U1411 ( .A(Dout[19]), .Y(aes_core_enc_block_n1400)
         );
  INVX1 aes_core_enc_block_U1410 ( .A(Dout[16]), .Y(aes_core_enc_block_n1426)
         );
  INVX1 aes_core_enc_block_U1409 ( .A(Dout[18]), .Y(aes_core_enc_block_n1448)
         );
  INVX1 aes_core_enc_block_U1408 ( .A(Dout[39]), .Y(aes_core_enc_block_n708)
         );
  INVX1 aes_core_enc_block_U1407 ( .A(Dout[28]), .Y(aes_core_enc_block_n1389)
         );
  INVX1 aes_core_enc_block_U1406 ( .A(Dout[25]), .Y(aes_core_enc_block_n1438)
         );
  INVX1 aes_core_enc_block_U1405 ( .A(Dout[43]), .Y(aes_core_enc_block_n1348)
         );
  INVX1 aes_core_enc_block_U1404 ( .A(Dout[42]), .Y(aes_core_enc_block_n189)
         );
  XNOR2X1 aes_core_enc_block_U1403 ( .A(aes_core_enc_block_n1420), .B(Dout[87]), .Y(aes_core_enc_block_n268) );
  XNOR2X1 aes_core_enc_block_U1402 ( .A(aes_core_enc_block_n1419), .B(Dout[63]), .Y(aes_core_enc_block_n741) );
  XNOR2X1 aes_core_enc_block_U1401 ( .A(aes_core_enc_block_n1416), .B(Dout[95]), .Y(aes_core_enc_block_n500) );
  XNOR2X1 aes_core_enc_block_U1400 ( .A(aes_core_enc_block_n1418), .B(Dout[31]), .Y(aes_core_enc_block_n980) );
  INVX1 aes_core_enc_block_U1399 ( .A(Dout[10]), .Y(aes_core_enc_block_n1458)
         );
  INVX1 aes_core_enc_block_U1398 ( .A(Dout[58]), .Y(aes_core_enc_block_n1441)
         );
  INVX1 aes_core_enc_block_U1397 ( .A(Dout[59]), .Y(aes_core_enc_block_n1453)
         );
  INVX1 aes_core_enc_block_U1396 ( .A(Dout[52]), .Y(aes_core_enc_block_n1401)
         );
  INVX1 aes_core_enc_block_U1395 ( .A(Dout[53]), .Y(aes_core_enc_block_n1406)
         );
  INVX1 aes_core_enc_block_U1394 ( .A(Dout[49]), .Y(aes_core_enc_block_n1431)
         );
  INVX1 aes_core_enc_block_U1393 ( .A(Dout[15]), .Y(aes_core_enc_block_n1371)
         );
  INVX1 aes_core_enc_block_U1392 ( .A(Dout[20]), .Y(aes_core_enc_block_n1390)
         );
  INVX1 aes_core_enc_block_U1391 ( .A(Dout[21]), .Y(aes_core_enc_block_n1405)
         );
  INVX1 aes_core_enc_block_U1390 ( .A(Dout[17]), .Y(aes_core_enc_block_n1439)
         );
  INVX1 aes_core_enc_block_U1389 ( .A(Dout[32]), .Y(aes_core_enc_block_n1396)
         );
  INVX1 aes_core_enc_block_U1388 ( .A(Dout[35]), .Y(aes_core_enc_block_n191)
         );
  INVX1 aes_core_enc_block_U1387 ( .A(Dout[34]), .Y(aes_core_enc_block_n1454)
         );
  INVX1 aes_core_enc_block_U1386 ( .A(Dout[63]), .Y(aes_core_enc_block_n1394)
         );
  INVX1 aes_core_enc_block_U1385 ( .A(Dout[0]), .Y(aes_core_enc_block_n947) );
  INVX1 aes_core_enc_block_U1384 ( .A(Dout[3]), .Y(aes_core_enc_block_n1455)
         );
  INVX1 aes_core_enc_block_U1383 ( .A(Dout[2]), .Y(aes_core_enc_block_n1457)
         );
  INVX1 aes_core_enc_block_U1382 ( .A(Dout[31]), .Y(aes_core_enc_block_n1383)
         );
  INVX1 aes_core_enc_block_U1381 ( .A(Dout[54]), .Y(aes_core_enc_block_n1412)
         );
  INVX1 aes_core_enc_block_U1380 ( .A(Dout[55]), .Y(aes_core_enc_block_n1416)
         );
  INVX1 aes_core_enc_block_U1379 ( .A(Dout[41]), .Y(aes_core_enc_block_n1363)
         );
  INVX1 aes_core_enc_block_U1378 ( .A(Dout[22]), .Y(aes_core_enc_block_n1411)
         );
  INVX1 aes_core_enc_block_U1377 ( .A(Dout[23]), .Y(aes_core_enc_block_n1419)
         );
  AOI221X1 aes_core_enc_block_U1376 ( .A0(aes_core_enc_block_n180), .A1(next), 
        .B0(aes_core_enc_block_n1185), .B1(aes_core_enc_block_n1195), .C0(
        aes_core_enc_block_n177), .Y(aes_core_enc_block_n1210) );
  INVX1 aes_core_enc_block_U1375 ( .A(aes_core_enc_block_n1210), .Y(
        aes_core_enc_block_n172) );
  INVX1 aes_core_enc_block_U1374 ( .A(Dout[60]), .Y(aes_core_enc_block_n1391)
         );
  INVX1 aes_core_enc_block_U1373 ( .A(Dout[61]), .Y(aes_core_enc_block_n1392)
         );
  INVX1 aes_core_enc_block_U1372 ( .A(Dout[62]), .Y(aes_core_enc_block_n1393)
         );
  INVX1 aes_core_enc_block_U1371 ( .A(Dout[57]), .Y(aes_core_enc_block_n1440)
         );
  INVX1 aes_core_enc_block_U1370 ( .A(Dout[5]), .Y(aes_core_enc_block_n195) );
  INVX1 aes_core_enc_block_U1369 ( .A(Dout[6]), .Y(aes_core_enc_block_n240) );
  INVX1 aes_core_enc_block_U1368 ( .A(Dout[4]), .Y(aes_core_enc_block_n192) );
  INVX1 aes_core_enc_block_U1367 ( .A(Dout[9]), .Y(aes_core_enc_block_n1373)
         );
  INVX1 aes_core_enc_block_U1366 ( .A(Dout[45]), .Y(aes_core_enc_block_n1353)
         );
  INVX1 aes_core_enc_block_U1365 ( .A(Dout[46]), .Y(aes_core_enc_block_n1356)
         );
  INVX1 aes_core_enc_block_U1364 ( .A(Dout[47]), .Y(aes_core_enc_block_n1359)
         );
  OAI32X1 aes_core_enc_block_U1363 ( .A0(aes_core_enc_block_n177), .A1(
        aes_core_enc_block_sword_ctr_reg[0]), .A2(aes_core_enc_block_n1209), 
        .B0(aes_core_enc_block_n173), .B1(aes_core_enc_block_n176), .Y(
        aes_core_enc_block_n1346) );
  XNOR2X1 aes_core_enc_block_U1362 ( .A(aes_core_enc_block_n1360), .B(Dout[15]), .Y(aes_core_enc_block_n619) );
  XNOR2X1 aes_core_enc_block_U1361 ( .A(aes_core_enc_block_n708), .B(Dout[79]), 
        .Y(aes_core_enc_block_n1099) );
  XNOR2X1 aes_core_enc_block_U1360 ( .A(aes_core_enc_block_n467), .B(Dout[71]), 
        .Y(aes_core_enc_block_n860) );
  XNOR2X1 aes_core_enc_block_U1359 ( .A(aes_core_enc_block_n1359), .B(Dout[7]), 
        .Y(aes_core_enc_block_n387) );
  INVX1 aes_core_enc_block_U1358 ( .A(Dout[36]), .Y(aes_core_enc_block_n1350)
         );
  INVX1 aes_core_enc_block_U1357 ( .A(Dout[37]), .Y(aes_core_enc_block_n194)
         );
  INVX1 aes_core_enc_block_U1356 ( .A(Dout[44]), .Y(aes_core_enc_block_n1377)
         );
  INVX1 aes_core_enc_block_U1355 ( .A(Dout[33]), .Y(aes_core_enc_block_n1456)
         );
  INVX1 aes_core_enc_block_U1354 ( .A(Dout[1]), .Y(aes_core_enc_block_n1397)
         );
  INVX1 aes_core_enc_block_U1353 ( .A(Dout[38]), .Y(aes_core_enc_block_n232)
         );
  INVX1 aes_core_enc_block_U1352 ( .A(Dout[8]), .Y(aes_core_enc_block_n1428)
         );
  XNOR2X1 aes_core_enc_block_U1351 ( .A(aes_core_enc_block_n1371), .B(Dout[55]), .Y(aes_core_enc_block_n476) );
  XNOR2X1 aes_core_enc_block_U1350 ( .A(aes_core_enc_block_n1359), .B(Dout[87]), .Y(aes_core_enc_block_n244) );
  XNOR2X1 aes_core_enc_block_U1349 ( .A(aes_core_enc_block_n467), .B(Dout[23]), 
        .Y(aes_core_enc_block_n717) );
  XNOR2X1 aes_core_enc_block_U1348 ( .A(aes_core_enc_block_n1418), .B(Dout[79]), .Y(aes_core_enc_block_n956) );
  AOI21X1 aes_core_enc_block_U1347 ( .A0(aes_core_enc_block_n180), .A1(
        aes_core_enc_block_enc_ctrl_reg[0]), .B0(aes_core_enc_block_n1194), 
        .Y(aes_core_enc_block_n1203) );
  XNOR2X1 aes_core_enc_block_U1346 ( .A(aes_core_enc_block_n1360), .B(Dout[95]), .Y(aes_core_enc_block_n542) );
  XNOR2X1 aes_core_enc_block_U1345 ( .A(aes_core_enc_block_n1383), .B(Dout[39]), .Y(aes_core_enc_block_n1022) );
  XNOR2X1 aes_core_enc_block_U1344 ( .A(aes_core_enc_block_n1394), .B(Dout[71]), .Y(aes_core_enc_block_n783) );
  XNOR2X1 aes_core_enc_block_U1343 ( .A(aes_core_enc_block_n1420), .B(Dout[7]), 
        .Y(aes_core_enc_block_n310) );
  XNOR2X1 aes_core_enc_block_U1342 ( .A(Dout[27]), .B(aes_core_enc_block_n972), 
        .Y(aes_core_enc_block_n1154) );
  XNOR2X1 aes_core_enc_block_U1341 ( .A(Dout[35]), .B(aes_core_enc_block_n1155), .Y(aes_core_enc_block_n1152) );
  XOR2X1 aes_core_enc_block_U1340 ( .A(aes_core_enc_block_n1154), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1153) );
  XOR2X1 aes_core_enc_block_U1339 ( .A(aes_core_enc_block_n1152), .B(
        aes_core_enc_block_n1153), .Y(aes_core_enc_block_n1151) );
  XNOR2X1 aes_core_enc_block_U1338 ( .A(Dout[0]), .B(aes_core_enc_block_n287), 
        .Y(aes_core_enc_block_n465) );
  XNOR2X1 aes_core_enc_block_U1337 ( .A(Dout[120]), .B(aes_core_enc_block_n466), .Y(aes_core_enc_block_n463) );
  XOR2X1 aes_core_enc_block_U1336 ( .A(aes_core_enc_block_n465), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n464) );
  XOR2X1 aes_core_enc_block_U1335 ( .A(aes_core_enc_block_n463), .B(
        aes_core_enc_block_n464), .Y(aes_core_enc_block_n462) );
  XNOR2X1 aes_core_enc_block_U1334 ( .A(Dout[12]), .B(aes_core_enc_block_n492), 
        .Y(aes_core_enc_block_n674) );
  XNOR2X1 aes_core_enc_block_U1333 ( .A(Dout[91]), .B(aes_core_enc_block_n675), 
        .Y(aes_core_enc_block_n672) );
  XOR2X1 aes_core_enc_block_U1332 ( .A(aes_core_enc_block_n674), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n673) );
  XOR2X1 aes_core_enc_block_U1331 ( .A(aes_core_enc_block_n672), .B(
        aes_core_enc_block_n673), .Y(aes_core_enc_block_n671) );
  XNOR2X1 aes_core_enc_block_U1330 ( .A(Dout[106]), .B(aes_core_enc_block_n717), .Y(aes_core_enc_block_n813) );
  XNOR2X1 aes_core_enc_block_U1329 ( .A(Dout[18]), .B(aes_core_enc_block_n814), 
        .Y(aes_core_enc_block_n811) );
  XOR2X1 aes_core_enc_block_U1328 ( .A(aes_core_enc_block_n813), .B(
        aes_core_enc_block_n750), .Y(aes_core_enc_block_n812) );
  XOR2X1 aes_core_enc_block_U1327 ( .A(aes_core_enc_block_n811), .B(
        aes_core_enc_block_n812), .Y(aes_core_enc_block_n810) );
  XNOR2X1 aes_core_enc_block_U1326 ( .A(Dout[11]), .B(aes_core_enc_block_n476), 
        .Y(aes_core_enc_block_n564) );
  XNOR2X1 aes_core_enc_block_U1325 ( .A(Dout[51]), .B(aes_core_enc_block_n565), 
        .Y(aes_core_enc_block_n562) );
  XOR2X1 aes_core_enc_block_U1324 ( .A(aes_core_enc_block_n564), .B(
        aes_core_enc_block_n501), .Y(aes_core_enc_block_n563) );
  XOR2X1 aes_core_enc_block_U1323 ( .A(aes_core_enc_block_n562), .B(
        aes_core_enc_block_n563), .Y(aes_core_enc_block_n561) );
  XNOR2X1 aes_core_enc_block_U1322 ( .A(Dout[123]), .B(aes_core_enc_block_n260), .Y(aes_core_enc_block_n442) );
  XNOR2X1 aes_core_enc_block_U1321 ( .A(Dout[3]), .B(aes_core_enc_block_n443), 
        .Y(aes_core_enc_block_n440) );
  XOR2X1 aes_core_enc_block_U1320 ( .A(aes_core_enc_block_n442), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n441) );
  XOR2X1 aes_core_enc_block_U1319 ( .A(aes_core_enc_block_n440), .B(
        aes_core_enc_block_n441), .Y(aes_core_enc_block_n439) );
  XNOR2X1 aes_core_enc_block_U1318 ( .A(Dout[11]), .B(aes_core_enc_block_n499), 
        .Y(aes_core_enc_block_n682) );
  XNOR2X1 aes_core_enc_block_U1317 ( .A(Dout[90]), .B(aes_core_enc_block_n683), 
        .Y(aes_core_enc_block_n680) );
  XOR2X1 aes_core_enc_block_U1316 ( .A(aes_core_enc_block_n682), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n681) );
  XOR2X1 aes_core_enc_block_U1315 ( .A(aes_core_enc_block_n680), .B(
        aes_core_enc_block_n681), .Y(aes_core_enc_block_n679) );
  XNOR2X1 aes_core_enc_block_U1314 ( .A(Dout[122]), .B(aes_core_enc_block_n267), .Y(aes_core_enc_block_n450) );
  XNOR2X1 aes_core_enc_block_U1313 ( .A(Dout[2]), .B(aes_core_enc_block_n451), 
        .Y(aes_core_enc_block_n448) );
  XOR2X1 aes_core_enc_block_U1312 ( .A(aes_core_enc_block_n450), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n449) );
  XOR2X1 aes_core_enc_block_U1311 ( .A(aes_core_enc_block_n448), .B(
        aes_core_enc_block_n449), .Y(aes_core_enc_block_n447) );
  XNOR2X1 aes_core_enc_block_U1310 ( .A(Dout[10]), .B(aes_core_enc_block_n476), 
        .Y(aes_core_enc_block_n572) );
  XNOR2X1 aes_core_enc_block_U1309 ( .A(Dout[50]), .B(aes_core_enc_block_n573), 
        .Y(aes_core_enc_block_n570) );
  XOR2X1 aes_core_enc_block_U1308 ( .A(aes_core_enc_block_n572), .B(
        aes_core_enc_block_n509), .Y(aes_core_enc_block_n571) );
  XOR2X1 aes_core_enc_block_U1307 ( .A(aes_core_enc_block_n570), .B(
        aes_core_enc_block_n571), .Y(aes_core_enc_block_n569) );
  XNOR2X1 aes_core_enc_block_U1306 ( .A(Dout[124]), .B(aes_core_enc_block_n244), .Y(aes_core_enc_block_n332) );
  XNOR2X1 aes_core_enc_block_U1305 ( .A(Dout[43]), .B(aes_core_enc_block_n333), 
        .Y(aes_core_enc_block_n330) );
  XOR2X1 aes_core_enc_block_U1304 ( .A(aes_core_enc_block_n332), .B(
        aes_core_enc_block_n269), .Y(aes_core_enc_block_n331) );
  XOR2X1 aes_core_enc_block_U1303 ( .A(aes_core_enc_block_n330), .B(
        aes_core_enc_block_n331), .Y(aes_core_enc_block_n329) );
  XNOR2X1 aes_core_enc_block_U1302 ( .A(Dout[115]), .B(aes_core_enc_block_n956), .Y(aes_core_enc_block_n1044) );
  XNOR2X1 aes_core_enc_block_U1301 ( .A(Dout[28]), .B(aes_core_enc_block_n1045), .Y(aes_core_enc_block_n1042) );
  XOR2X1 aes_core_enc_block_U1300 ( .A(aes_core_enc_block_n1044), .B(
        aes_core_enc_block_n981), .Y(aes_core_enc_block_n1043) );
  XOR2X1 aes_core_enc_block_U1299 ( .A(aes_core_enc_block_n1042), .B(
        aes_core_enc_block_n1043), .Y(aes_core_enc_block_n1041) );
  XNOR2X1 aes_core_enc_block_U1298 ( .A(Dout[114]), .B(aes_core_enc_block_n956), .Y(aes_core_enc_block_n1052) );
  XNOR2X1 aes_core_enc_block_U1297 ( .A(Dout[27]), .B(aes_core_enc_block_n1053), .Y(aes_core_enc_block_n1050) );
  XOR2X1 aes_core_enc_block_U1296 ( .A(aes_core_enc_block_n1052), .B(
        aes_core_enc_block_n989), .Y(aes_core_enc_block_n1051) );
  XOR2X1 aes_core_enc_block_U1295 ( .A(aes_core_enc_block_n1050), .B(
        aes_core_enc_block_n1051), .Y(aes_core_enc_block_n1049) );
  XNOR2X1 aes_core_enc_block_U1294 ( .A(Dout[107]), .B(aes_core_enc_block_n717), .Y(aes_core_enc_block_n805) );
  XNOR2X1 aes_core_enc_block_U1293 ( .A(Dout[19]), .B(aes_core_enc_block_n806), 
        .Y(aes_core_enc_block_n803) );
  XOR2X1 aes_core_enc_block_U1292 ( .A(aes_core_enc_block_n805), .B(
        aes_core_enc_block_n742), .Y(aes_core_enc_block_n804) );
  XOR2X1 aes_core_enc_block_U1291 ( .A(aes_core_enc_block_n803), .B(
        aes_core_enc_block_n804), .Y(aes_core_enc_block_n802) );
  XNOR2X1 aes_core_enc_block_U1290 ( .A(Dout[121]), .B(aes_core_enc_block_n244), .Y(aes_core_enc_block_n355) );
  XNOR2X1 aes_core_enc_block_U1289 ( .A(Dout[40]), .B(aes_core_enc_block_n356), 
        .Y(aes_core_enc_block_n353) );
  XOR2X1 aes_core_enc_block_U1288 ( .A(aes_core_enc_block_n355), .B(
        aes_core_enc_block_n294), .Y(aes_core_enc_block_n354) );
  XOR2X1 aes_core_enc_block_U1287 ( .A(aes_core_enc_block_n353), .B(
        aes_core_enc_block_n354), .Y(aes_core_enc_block_n352) );
  XNOR2X1 aes_core_enc_block_U1286 ( .A(Dout[123]), .B(aes_core_enc_block_n244), .Y(aes_core_enc_block_n340) );
  XNOR2X1 aes_core_enc_block_U1285 ( .A(Dout[42]), .B(aes_core_enc_block_n341), 
        .Y(aes_core_enc_block_n338) );
  XOR2X1 aes_core_enc_block_U1284 ( .A(aes_core_enc_block_n340), .B(
        aes_core_enc_block_n277), .Y(aes_core_enc_block_n339) );
  XOR2X1 aes_core_enc_block_U1283 ( .A(aes_core_enc_block_n338), .B(
        aes_core_enc_block_n339), .Y(aes_core_enc_block_n337) );
  XNOR2X1 aes_core_enc_block_U1282 ( .A(Dout[26]), .B(aes_core_enc_block_n979), 
        .Y(aes_core_enc_block_n1162) );
  XNOR2X1 aes_core_enc_block_U1281 ( .A(Dout[34]), .B(aes_core_enc_block_n1163), .Y(aes_core_enc_block_n1160) );
  XOR2X1 aes_core_enc_block_U1280 ( .A(aes_core_enc_block_n1162), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1161) );
  XOR2X1 aes_core_enc_block_U1279 ( .A(aes_core_enc_block_n1160), .B(
        aes_core_enc_block_n1161), .Y(aes_core_enc_block_n1159) );
  XNOR2X1 aes_core_enc_block_U1278 ( .A(aes_core_enc_block_n140), .B(Dout[103]), .Y(aes_core_enc_block_n473) );
  XNOR2X1 aes_core_enc_block_U1277 ( .A(aes_core_enc_block_n166), .B(Dout[117]), .Y(aes_core_enc_block_n969) );
  XNOR2X1 aes_core_enc_block_U1276 ( .A(aes_core_enc_block_n165), .B(Dout[118]), .Y(aes_core_enc_block_n961) );
  XNOR2X1 aes_core_enc_block_U1275 ( .A(aes_core_enc_block_n171), .B(Dout[112]), .Y(aes_core_enc_block_n1013) );
  XNOR2X1 aes_core_enc_block_U1274 ( .A(aes_core_enc_block_n169), .B(Dout[114]), .Y(aes_core_enc_block_n996) );
  XNOR2X1 aes_core_enc_block_U1273 ( .A(aes_core_enc_block_n142), .B(Dout[53]), 
        .Y(aes_core_enc_block_n489) );
  XNOR2X1 aes_core_enc_block_U1272 ( .A(aes_core_enc_block_n141), .B(Dout[54]), 
        .Y(aes_core_enc_block_n481) );
  XNOR2X1 aes_core_enc_block_U1271 ( .A(aes_core_enc_block_n150), .B(Dout[21]), 
        .Y(aes_core_enc_block_n730) );
  XNOR2X1 aes_core_enc_block_U1270 ( .A(aes_core_enc_block_n149), .B(Dout[22]), 
        .Y(aes_core_enc_block_n722) );
  XNOR2X1 aes_core_enc_block_U1269 ( .A(aes_core_enc_block_n135), .B(Dout[84]), 
        .Y(aes_core_enc_block_n270) );
  XOR2X1 aes_core_enc_block_U1268 ( .A(aes_core_enc_block_n269), .B(
        aes_core_enc_block_n270), .Y(aes_core_enc_block_n265) );
  XNOR2X1 aes_core_enc_block_U1267 ( .A(aes_core_enc_block_n167), .B(Dout[116]), .Y(aes_core_enc_block_n982) );
  XOR2X1 aes_core_enc_block_U1266 ( .A(aes_core_enc_block_n981), .B(
        aes_core_enc_block_n982), .Y(aes_core_enc_block_n977) );
  XNOR2X1 aes_core_enc_block_U1265 ( .A(aes_core_enc_block_n151), .B(Dout[20]), 
        .Y(aes_core_enc_block_n743) );
  XOR2X1 aes_core_enc_block_U1264 ( .A(aes_core_enc_block_n742), .B(
        aes_core_enc_block_n743), .Y(aes_core_enc_block_n738) );
  XNOR2X1 aes_core_enc_block_U1263 ( .A(aes_core_enc_block_n143), .B(Dout[52]), 
        .Y(aes_core_enc_block_n502) );
  XOR2X1 aes_core_enc_block_U1262 ( .A(aes_core_enc_block_n501), .B(
        aes_core_enc_block_n502), .Y(aes_core_enc_block_n497) );
  XNOR2X1 aes_core_enc_block_U1261 ( .A(aes_core_enc_block_n134), .B(Dout[85]), 
        .Y(aes_core_enc_block_n257) );
  XNOR2X1 aes_core_enc_block_U1260 ( .A(aes_core_enc_block_n133), .B(Dout[86]), 
        .Y(aes_core_enc_block_n249) );
  XNOR2X1 aes_core_enc_block_U1259 ( .A(aes_core_enc_block_n139), .B(Dout[80]), 
        .Y(aes_core_enc_block_n301) );
  XNOR2X1 aes_core_enc_block_U1258 ( .A(aes_core_enc_block_n137), .B(Dout[82]), 
        .Y(aes_core_enc_block_n284) );
  XNOR2X1 aes_core_enc_block_U1257 ( .A(aes_core_enc_block_n147), .B(Dout[48]), 
        .Y(aes_core_enc_block_n533) );
  XNOR2X1 aes_core_enc_block_U1256 ( .A(aes_core_enc_block_n145), .B(Dout[50]), 
        .Y(aes_core_enc_block_n516) );
  XNOR2X1 aes_core_enc_block_U1255 ( .A(aes_core_enc_block_n155), .B(Dout[16]), 
        .Y(aes_core_enc_block_n774) );
  XNOR2X1 aes_core_enc_block_U1254 ( .A(aes_core_enc_block_n153), .B(Dout[18]), 
        .Y(aes_core_enc_block_n757) );
  XNOR2X1 aes_core_enc_block_U1253 ( .A(aes_core_enc_block_n156), .B(Dout[39]), 
        .Y(aes_core_enc_block_n953) );
  XNOR2X1 aes_core_enc_block_U1252 ( .A(aes_core_enc_block_n146), .B(Dout[49]), 
        .Y(aes_core_enc_block_n528) );
  XOR2X1 aes_core_enc_block_U1251 ( .A(aes_core_enc_block_n500), .B(
        aes_core_enc_block_n528), .Y(aes_core_enc_block_n524) );
  XNOR2X1 aes_core_enc_block_U1250 ( .A(aes_core_enc_block_n138), .B(Dout[81]), 
        .Y(aes_core_enc_block_n296) );
  XOR2X1 aes_core_enc_block_U1249 ( .A(aes_core_enc_block_n268), .B(
        aes_core_enc_block_n296), .Y(aes_core_enc_block_n292) );
  XNOR2X1 aes_core_enc_block_U1248 ( .A(aes_core_enc_block_n170), .B(Dout[113]), .Y(aes_core_enc_block_n1008) );
  XOR2X1 aes_core_enc_block_U1247 ( .A(aes_core_enc_block_n980), .B(
        aes_core_enc_block_n1008), .Y(aes_core_enc_block_n1004) );
  XNOR2X1 aes_core_enc_block_U1246 ( .A(aes_core_enc_block_n154), .B(Dout[17]), 
        .Y(aes_core_enc_block_n769) );
  XOR2X1 aes_core_enc_block_U1245 ( .A(aes_core_enc_block_n741), .B(
        aes_core_enc_block_n769), .Y(aes_core_enc_block_n765) );
  XNOR2X1 aes_core_enc_block_U1244 ( .A(aes_core_enc_block_n136), .B(Dout[83]), 
        .Y(aes_core_enc_block_n279) );
  XOR2X1 aes_core_enc_block_U1243 ( .A(aes_core_enc_block_n268), .B(
        aes_core_enc_block_n279), .Y(aes_core_enc_block_n275) );
  XNOR2X1 aes_core_enc_block_U1242 ( .A(aes_core_enc_block_n168), .B(Dout[115]), .Y(aes_core_enc_block_n991) );
  XOR2X1 aes_core_enc_block_U1241 ( .A(aes_core_enc_block_n980), .B(
        aes_core_enc_block_n991), .Y(aes_core_enc_block_n987) );
  XNOR2X1 aes_core_enc_block_U1240 ( .A(aes_core_enc_block_n144), .B(Dout[51]), 
        .Y(aes_core_enc_block_n511) );
  XOR2X1 aes_core_enc_block_U1239 ( .A(aes_core_enc_block_n500), .B(
        aes_core_enc_block_n511), .Y(aes_core_enc_block_n507) );
  XNOR2X1 aes_core_enc_block_U1238 ( .A(aes_core_enc_block_n152), .B(Dout[19]), 
        .Y(aes_core_enc_block_n752) );
  XOR2X1 aes_core_enc_block_U1237 ( .A(aes_core_enc_block_n741), .B(
        aes_core_enc_block_n752), .Y(aes_core_enc_block_n748) );
  XNOR2X1 aes_core_enc_block_U1236 ( .A(aes_core_enc_block_n148), .B(Dout[71]), 
        .Y(aes_core_enc_block_n714) );
  XNOR2X1 aes_core_enc_block_U1235 ( .A(Dout[24]), .B(aes_core_enc_block_n999), 
        .Y(aes_core_enc_block_n1177) );
  XNOR2X1 aes_core_enc_block_U1234 ( .A(Dout[32]), .B(aes_core_enc_block_n1178), .Y(aes_core_enc_block_n1175) );
  XOR2X1 aes_core_enc_block_U1233 ( .A(aes_core_enc_block_n1177), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1176) );
  XOR2X1 aes_core_enc_block_U1232 ( .A(aes_core_enc_block_n1175), .B(
        aes_core_enc_block_n1176), .Y(aes_core_enc_block_n1174) );
  XNOR2X1 aes_core_enc_block_U1231 ( .A(Dout[88]), .B(aes_core_enc_block_n519), 
        .Y(aes_core_enc_block_n697) );
  XNOR2X1 aes_core_enc_block_U1230 ( .A(Dout[96]), .B(aes_core_enc_block_n698), 
        .Y(aes_core_enc_block_n695) );
  XOR2X1 aes_core_enc_block_U1229 ( .A(aes_core_enc_block_n697), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n696) );
  XOR2X1 aes_core_enc_block_U1228 ( .A(aes_core_enc_block_n695), .B(
        aes_core_enc_block_n696), .Y(aes_core_enc_block_n694) );
  XNOR2X1 aes_core_enc_block_U1227 ( .A(aes_core_enc_block_n132), .B(Dout[7]), 
        .Y(aes_core_enc_block_n241) );
  XNOR2X1 aes_core_enc_block_U1226 ( .A(Dout[104]), .B(aes_core_enc_block_n717), .Y(aes_core_enc_block_n828) );
  XNOR2X1 aes_core_enc_block_U1225 ( .A(Dout[16]), .B(aes_core_enc_block_n829), 
        .Y(aes_core_enc_block_n826) );
  XOR2X1 aes_core_enc_block_U1224 ( .A(aes_core_enc_block_n828), .B(
        aes_core_enc_block_n767), .Y(aes_core_enc_block_n827) );
  XOR2X1 aes_core_enc_block_U1223 ( .A(aes_core_enc_block_n826), .B(
        aes_core_enc_block_n827), .Y(aes_core_enc_block_n825) );
  XNOR2X1 aes_core_enc_block_U1222 ( .A(Dout[48]), .B(aes_core_enc_block_n476), 
        .Y(aes_core_enc_block_n587) );
  XNOR2X1 aes_core_enc_block_U1221 ( .A(Dout[89]), .B(aes_core_enc_block_n588), 
        .Y(aes_core_enc_block_n585) );
  XOR2X1 aes_core_enc_block_U1220 ( .A(aes_core_enc_block_n587), .B(
        aes_core_enc_block_n526), .Y(aes_core_enc_block_n586) );
  XOR2X1 aes_core_enc_block_U1219 ( .A(aes_core_enc_block_n585), .B(
        aes_core_enc_block_n586), .Y(aes_core_enc_block_n584) );
  XNOR2X1 aes_core_enc_block_U1218 ( .A(Dout[107]), .B(aes_core_enc_block_n740), .Y(aes_core_enc_block_n923) );
  XNOR2X1 aes_core_enc_block_U1217 ( .A(Dout[58]), .B(aes_core_enc_block_n924), 
        .Y(aes_core_enc_block_n921) );
  XOR2X1 aes_core_enc_block_U1216 ( .A(aes_core_enc_block_n923), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n922) );
  XOR2X1 aes_core_enc_block_U1215 ( .A(aes_core_enc_block_n921), .B(
        aes_core_enc_block_n922), .Y(aes_core_enc_block_n920) );
  XNOR2X1 aes_core_enc_block_U1214 ( .A(Dout[108]), .B(aes_core_enc_block_n733), .Y(aes_core_enc_block_n915) );
  XNOR2X1 aes_core_enc_block_U1213 ( .A(Dout[59]), .B(aes_core_enc_block_n916), 
        .Y(aes_core_enc_block_n913) );
  XOR2X1 aes_core_enc_block_U1212 ( .A(aes_core_enc_block_n915), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n914) );
  XOR2X1 aes_core_enc_block_U1211 ( .A(aes_core_enc_block_n913), .B(
        aes_core_enc_block_n914), .Y(aes_core_enc_block_n912) );
  XNOR2X1 aes_core_enc_block_U1210 ( .A(Dout[105]), .B(aes_core_enc_block_n760), .Y(aes_core_enc_block_n938) );
  XNOR2X1 aes_core_enc_block_U1209 ( .A(Dout[56]), .B(aes_core_enc_block_n939), 
        .Y(aes_core_enc_block_n936) );
  XOR2X1 aes_core_enc_block_U1208 ( .A(aes_core_enc_block_n938), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n937) );
  XOR2X1 aes_core_enc_block_U1207 ( .A(aes_core_enc_block_n936), .B(
        aes_core_enc_block_n937), .Y(aes_core_enc_block_n935) );
  XNOR2X1 aes_core_enc_block_U1206 ( .A(Dout[112]), .B(aes_core_enc_block_n956), .Y(aes_core_enc_block_n1067) );
  XNOR2X1 aes_core_enc_block_U1205 ( .A(Dout[25]), .B(aes_core_enc_block_n1068), .Y(aes_core_enc_block_n1065) );
  XOR2X1 aes_core_enc_block_U1204 ( .A(aes_core_enc_block_n1067), .B(
        aes_core_enc_block_n1006), .Y(aes_core_enc_block_n1066) );
  XOR2X1 aes_core_enc_block_U1203 ( .A(aes_core_enc_block_n1065), .B(
        aes_core_enc_block_n1066), .Y(aes_core_enc_block_n1064) );
  OAI22X1 aes_core_enc_block_U1202 ( .A0(Din[125]), .A1(aes_core_enc_block_n99), .B0(Dout[125]), .B1(aes_core_enc_block_n26), .Y(aes_core_enc_block_n256) );
  OAI22X1 aes_core_enc_block_U1201 ( .A0(Din[126]), .A1(aes_core_enc_block_n99), .B0(Dout[126]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n248) );
  OAI22X1 aes_core_enc_block_U1200 ( .A0(Din[127]), .A1(aes_core_enc_block_n99), .B0(Dout[127]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n238) );
  OAI22X1 aes_core_enc_block_U1199 ( .A0(Din[124]), .A1(aes_core_enc_block_n99), .B0(Dout[124]), .B1(aes_core_enc_block_n26), .Y(aes_core_enc_block_n264) );
  OAI22X1 aes_core_enc_block_U1198 ( .A0(Din[120]), .A1(aes_core_enc_block_n99), .B0(Dout[120]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n300) );
  OAI22X1 aes_core_enc_block_U1197 ( .A0(Din[121]), .A1(aes_core_enc_block_n99), .B0(Dout[121]), .B1(aes_core_enc_block_n26), .Y(aes_core_enc_block_n291) );
  OAI22X1 aes_core_enc_block_U1196 ( .A0(Din[122]), .A1(aes_core_enc_block_n99), .B0(Dout[122]), .B1(aes_core_enc_block_n26), .Y(aes_core_enc_block_n283) );
  OAI22X1 aes_core_enc_block_U1195 ( .A0(Din[92]), .A1(aes_core_enc_block_n99), 
        .B0(Dout[92]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n496) );
  OAI22X1 aes_core_enc_block_U1194 ( .A0(Din[93]), .A1(aes_core_enc_block_n94), 
        .B0(Dout[93]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n488) );
  OAI22X1 aes_core_enc_block_U1193 ( .A0(Din[94]), .A1(aes_core_enc_block_n99), 
        .B0(Dout[94]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n480) );
  OAI22X1 aes_core_enc_block_U1192 ( .A0(Din[123]), .A1(aes_core_enc_block_n99), .B0(Dout[123]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n274) );
  OAI22X1 aes_core_enc_block_U1191 ( .A0(Din[88]), .A1(aes_core_enc_block_n100), .B0(Dout[88]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n532) );
  OAI22X1 aes_core_enc_block_U1190 ( .A0(Din[89]), .A1(aes_core_enc_block_n95), 
        .B0(Dout[89]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n523) );
  OAI22X1 aes_core_enc_block_U1189 ( .A0(Din[90]), .A1(aes_core_enc_block_n100), .B0(Dout[90]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n515) );
  OAI22X1 aes_core_enc_block_U1188 ( .A0(Din[91]), .A1(aes_core_enc_block_n95), 
        .B0(Dout[91]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n506) );
  OAI22X1 aes_core_enc_block_U1187 ( .A0(Din[60]), .A1(aes_core_enc_block_n100), .B0(Dout[60]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n737) );
  OAI22X1 aes_core_enc_block_U1186 ( .A0(Din[61]), .A1(aes_core_enc_block_n95), 
        .B0(Dout[61]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n729) );
  OAI22X1 aes_core_enc_block_U1185 ( .A0(Din[62]), .A1(aes_core_enc_block_n100), .B0(Dout[62]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n721) );
  OAI22X1 aes_core_enc_block_U1184 ( .A0(Din[63]), .A1(aes_core_enc_block_n94), 
        .B0(Dout[63]), .B1(aes_core_enc_block_n27), .Y(aes_core_enc_block_n713) );
  OAI22X1 aes_core_enc_block_U1183 ( .A0(Din[57]), .A1(aes_core_enc_block_n95), 
        .B0(Dout[57]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n764) );
  OAI22X1 aes_core_enc_block_U1182 ( .A0(Din[29]), .A1(aes_core_enc_block_n100), .B0(Dout[29]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n968) );
  OAI22X1 aes_core_enc_block_U1181 ( .A0(Din[30]), .A1(aes_core_enc_block_n100), .B0(Dout[30]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n960) );
  OAI22X1 aes_core_enc_block_U1180 ( .A0(Din[31]), .A1(aes_core_enc_block_n100), .B0(Dout[31]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n952) );
  OAI22X1 aes_core_enc_block_U1179 ( .A0(Din[95]), .A1(aes_core_enc_block_n94), 
        .B0(Dout[95]), .B1(aes_core_enc_block_n26), .Y(aes_core_enc_block_n472) );
  OAI22X1 aes_core_enc_block_U1178 ( .A0(Din[56]), .A1(aes_core_enc_block_n99), 
        .B0(Dout[56]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n773) );
  OAI22X1 aes_core_enc_block_U1177 ( .A0(Din[58]), .A1(aes_core_enc_block_n100), .B0(Dout[58]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n756) );
  OAI22X1 aes_core_enc_block_U1176 ( .A0(Din[59]), .A1(aes_core_enc_block_n95), 
        .B0(Dout[59]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n747) );
  OAI22X1 aes_core_enc_block_U1175 ( .A0(Din[28]), .A1(aes_core_enc_block_n99), 
        .B0(Dout[28]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n976) );
  OAI22X1 aes_core_enc_block_U1174 ( .A0(Din[24]), .A1(aes_core_enc_block_n100), .B0(Dout[24]), .B1(aes_core_enc_block_n76), .Y(aes_core_enc_block_n1012) );
  OAI22X1 aes_core_enc_block_U1173 ( .A0(Din[25]), .A1(aes_core_enc_block_n100), .B0(Dout[25]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n1003) );
  OAI22X1 aes_core_enc_block_U1172 ( .A0(Din[26]), .A1(aes_core_enc_block_n100), .B0(Dout[26]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n995) );
  OAI22X1 aes_core_enc_block_U1171 ( .A0(Din[27]), .A1(aes_core_enc_block_n100), .B0(Dout[27]), .B1(aes_core_enc_block_n28), .Y(aes_core_enc_block_n986) );
  INVX1 aes_core_enc_block_U1170 ( .A(Dout[71]), .Y(aes_core_enc_block_n1415)
         );
  INVX1 aes_core_enc_block_U1169 ( .A(Dout[79]), .Y(aes_core_enc_block_n1382)
         );
  INVX1 aes_core_enc_block_U1168 ( .A(Dout[87]), .Y(aes_core_enc_block_n1417)
         );
  INVX1 aes_core_enc_block_U1167 ( .A(Dout[95]), .Y(aes_core_enc_block_n1361)
         );
  INVX1 aes_core_enc_block_U1166 ( .A(Dout[103]), .Y(aes_core_enc_block_n1360)
         );
  INVX1 aes_core_enc_block_U1165 ( .A(Dout[126]), .Y(aes_core_enc_block_n1409)
         );
  INVX1 aes_core_enc_block_U1164 ( .A(Dout[127]), .Y(aes_core_enc_block_n1420)
         );
  INVX1 aes_core_enc_block_U1163 ( .A(Dout[111]), .Y(aes_core_enc_block_n467)
         );
  INVX1 aes_core_enc_block_U1162 ( .A(Dout[119]), .Y(aes_core_enc_block_n1418)
         );
  INVX1 aes_core_enc_block_U1161 ( .A(Dout[86]), .Y(aes_core_enc_block_n1414)
         );
  INVX1 aes_core_enc_block_U1160 ( .A(Dout[118]), .Y(aes_core_enc_block_n1410)
         );
  INVX1 aes_core_enc_block_U1159 ( .A(Dout[78]), .Y(aes_core_enc_block_n1370)
         );
  INVX1 aes_core_enc_block_U1158 ( .A(Dout[94]), .Y(aes_core_enc_block_n1413)
         );
  INVX1 aes_core_enc_block_U1157 ( .A(Dout[70]), .Y(aes_core_enc_block_n1358)
         );
  INVX1 aes_core_enc_block_U1156 ( .A(Dout[110]), .Y(aes_core_enc_block_n196)
         );
  INVX1 aes_core_enc_block_U1155 ( .A(Dout[102]), .Y(aes_core_enc_block_n1357)
         );
  INVX1 aes_core_enc_block_U1154 ( .A(Dout[114]), .Y(aes_core_enc_block_n1446)
         );
  INVX1 aes_core_enc_block_U1153 ( .A(Dout[90]), .Y(aes_core_enc_block_n1443)
         );
  INVX1 aes_core_enc_block_U1152 ( .A(Dout[85]), .Y(aes_core_enc_block_n1407)
         );
  INVX1 aes_core_enc_block_U1151 ( .A(Dout[82]), .Y(aes_core_enc_block_n1444)
         );
  INVX1 aes_core_enc_block_U1150 ( .A(Dout[106]), .Y(aes_core_enc_block_n1364)
         );
  INVX1 aes_core_enc_block_U1149 ( .A(Dout[117]), .Y(aes_core_enc_block_n1378)
         );
  INVX1 aes_core_enc_block_U1148 ( .A(Dout[122]), .Y(aes_core_enc_block_n1445)
         );
  INVX1 aes_core_enc_block_U1147 ( .A(Dout[98]), .Y(aes_core_enc_block_n1398)
         );
  INVX1 aes_core_enc_block_U1146 ( .A(Dout[69]), .Y(aes_core_enc_block_n1355)
         );
  INVX1 aes_core_enc_block_U1145 ( .A(Dout[66]), .Y(aes_core_enc_block_n1347)
         );
  INVX1 aes_core_enc_block_U1144 ( .A(Dout[74]), .Y(aes_core_enc_block_n1374)
         );
  INVX1 aes_core_enc_block_U1143 ( .A(Dout[93]), .Y(aes_core_enc_block_n1403)
         );
  INVX1 aes_core_enc_block_U1142 ( .A(Dout[125]), .Y(aes_core_enc_block_n1408)
         );
  INVX1 aes_core_enc_block_U1141 ( .A(Dout[101]), .Y(aes_core_enc_block_n1354)
         );
  OAI221X1 aes_core_enc_block_U1140 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1361), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1420), .C0(aes_core_enc_block_n205), .Y(
        aes_core_enc_sboxw[31]) );
  AOI22X1 aes_core_enc_block_U1139 ( .A0(Dout[31]), .A1(aes_core_enc_block_n11), .B0(Dout[63]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n205) );
  INVX1 aes_core_enc_block_U1138 ( .A(Dout[107]), .Y(aes_core_enc_block_n190)
         );
  INVX1 aes_core_enc_block_U1137 ( .A(Dout[115]), .Y(aes_core_enc_block_n1450)
         );
  INVX1 aes_core_enc_block_U1136 ( .A(Dout[112]), .Y(aes_core_enc_block_n1424)
         );
  INVX1 aes_core_enc_block_U1135 ( .A(Dout[123]), .Y(aes_core_enc_block_n1449)
         );
  INVX1 aes_core_enc_block_U1134 ( .A(Dout[89]), .Y(aes_core_enc_block_n1432)
         );
  INVX1 aes_core_enc_block_U1133 ( .A(Dout[96]), .Y(aes_core_enc_block_n187)
         );
  INVX1 aes_core_enc_block_U1132 ( .A(Dout[84]), .Y(aes_core_enc_block_n1366)
         );
  INVX1 aes_core_enc_block_U1131 ( .A(Dout[80]), .Y(aes_core_enc_block_n1430)
         );
  INVX1 aes_core_enc_block_U1130 ( .A(Dout[81]), .Y(aes_core_enc_block_n1433)
         );
  INVX1 aes_core_enc_block_U1129 ( .A(Dout[83]), .Y(aes_core_enc_block_n1386)
         );
  INVX1 aes_core_enc_block_U1128 ( .A(Dout[88]), .Y(aes_core_enc_block_n1429)
         );
  INVX1 aes_core_enc_block_U1127 ( .A(Dout[91]), .Y(aes_core_enc_block_n1452)
         );
  INVX1 aes_core_enc_block_U1126 ( .A(Dout[105]), .Y(aes_core_enc_block_n1436)
         );
  INVX1 aes_core_enc_block_U1125 ( .A(Dout[108]), .Y(aes_core_enc_block_n1349)
         );
  INVX1 aes_core_enc_block_U1124 ( .A(Dout[116]), .Y(aes_core_enc_block_n1388)
         );
  INVX1 aes_core_enc_block_U1123 ( .A(Dout[113]), .Y(aes_core_enc_block_n1435)
         );
  INVX1 aes_core_enc_block_U1122 ( .A(Dout[124]), .Y(aes_core_enc_block_n1387)
         );
  INVX1 aes_core_enc_block_U1121 ( .A(Dout[121]), .Y(aes_core_enc_block_n1434)
         );
  INVX1 aes_core_enc_block_U1120 ( .A(Dout[104]), .Y(aes_core_enc_block_n1422)
         );
  INVX1 aes_core_enc_block_U1119 ( .A(Dout[120]), .Y(aes_core_enc_block_n1421)
         );
  INVX1 aes_core_enc_block_U1118 ( .A(Dout[99]), .Y(aes_core_enc_block_n1385)
         );
  INVX1 aes_core_enc_block_U1117 ( .A(Dout[67]), .Y(aes_core_enc_block_n1376)
         );
  INVX1 aes_core_enc_block_U1116 ( .A(Dout[68]), .Y(aes_core_enc_block_n1352)
         );
  INVX1 aes_core_enc_block_U1115 ( .A(Dout[76]), .Y(aes_core_enc_block_n1368)
         );
  INVX1 aes_core_enc_block_U1114 ( .A(Dout[77]), .Y(aes_core_enc_block_n1404)
         );
  INVX1 aes_core_enc_block_U1113 ( .A(Dout[73]), .Y(aes_core_enc_block_n1437)
         );
  INVX1 aes_core_enc_block_U1112 ( .A(Dout[75]), .Y(aes_core_enc_block_n1399)
         );
  INVX1 aes_core_enc_block_U1110 ( .A(Dout[72]), .Y(aes_core_enc_block_n1372)
         );
  INVX1 aes_core_enc_block_U1109 ( .A(Dout[65]), .Y(aes_core_enc_block_n188)
         );
  INVX1 aes_core_enc_block_U1108 ( .A(Dout[92]), .Y(aes_core_enc_block_n1402)
         );
  INVX1 aes_core_enc_block_U1107 ( .A(Dout[109]), .Y(aes_core_enc_block_n193)
         );
  INVX1 aes_core_enc_block_U1106 ( .A(Dout[100]), .Y(aes_core_enc_block_n1367)
         );
  INVX1 aes_core_enc_block_U1105 ( .A(Dout[97]), .Y(aes_core_enc_block_n1207)
         );
  OAI221X1 aes_core_enc_block_U1104 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1417), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1418), .C0(aes_core_enc_block_n214), .Y(
        aes_core_enc_sboxw[23]) );
  OAI221X1 aes_core_enc_block_U1103 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1414), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1410), .C0(aes_core_enc_block_n215), .Y(
        aes_core_enc_sboxw[22]) );
  OAI221X1 aes_core_enc_block_U1102 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1382), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n467), .C0(aes_core_enc_block_n223), .Y(
        aes_core_enc_sboxw[15]) );
  OAI221X1 aes_core_enc_block_U1101 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1415), .B0(aes_core_enc_block_n127), .B1(
        aes_core_enc_block_n1360), .C0(aes_core_enc_block_n200), .Y(
        aes_core_enc_sboxw[7]) );
  OAI221X1 aes_core_enc_block_U1100 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1370), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n196), .C0(aes_core_enc_block_n224), .Y(
        aes_core_enc_sboxw[14]) );
  OAI221X1 aes_core_enc_block_U1099 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1358), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1357), .C0(aes_core_enc_block_n201), .Y(
        aes_core_enc_sboxw[6]) );
  OAI221X1 aes_core_enc_block_U1098 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1413), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1409), .C0(aes_core_enc_block_n206), .Y(
        aes_core_enc_sboxw[30]) );
  AOI22X1 aes_core_enc_block_U1097 ( .A0(Dout[6]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[38]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n201) );
  AOI22X1 aes_core_enc_block_U1096 ( .A0(Dout[14]), .A1(aes_core_enc_block_n10), .B0(Dout[46]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n224) );
  AOI22X1 aes_core_enc_block_U1095 ( .A0(Dout[15]), .A1(aes_core_enc_block_n10), .B0(Dout[47]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n223) );
  AOI22X1 aes_core_enc_block_U1094 ( .A0(Dout[23]), .A1(aes_core_enc_block_n10), .B0(Dout[55]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n214) );
  AOI22X1 aes_core_enc_block_U1093 ( .A0(Dout[22]), .A1(aes_core_enc_block_n10), .B0(Dout[54]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n215) );
  AOI22X1 aes_core_enc_block_U1092 ( .A0(Dout[30]), .A1(aes_core_enc_block_n10), .B0(Dout[62]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n206) );
  AOI22X1 aes_core_enc_block_U1091 ( .A0(Dout[7]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[39]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n200) );
  NOR2X1 aes_core_enc_block_U1090 ( .A(aes_core_enc_block_n174), .B(
        aes_core_enc_block_sword_ctr_reg[0]), .Y(aes_core_enc_block_n946) );
  NOR2X1 aes_core_enc_block_U1089 ( .A(aes_core_enc_block_n173), .B(
        aes_core_enc_block_sword_ctr_reg[1]), .Y(aes_core_enc_block_n707) );
  XOR2X1 aes_core_enc_block_U1088 ( .A(aes_core_enc_block_n987), .B(
        aes_core_enc_block_n988), .Y(aes_core_enc_block_n984) );
  OAI2BB2X1 aes_core_enc_block_U1087 ( .B0(aes_core_enc_block_n1451), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n116), .A1N(Din[27]), 
        .Y(aes_core_enc_block_n985) );
  AOI222X1 aes_core_enc_block_U1086 ( .A0(aes_core_enc_block_n118), .A1(
        aes_core_enc_block_n984), .B0(aes_core_enc_block_n985), .B1(
        aes_core_enc_block_n168), .C0(aes_core_round_key[27]), .C1(
        aes_core_enc_block_n986), .Y(aes_core_enc_block_n983) );
  OAI221X1 aes_core_enc_block_U1085 ( .A0(aes_core_enc_block_n162), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1451), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n983), .Y(
        aes_core_enc_block_n1310) );
  XNOR2X1 aes_core_enc_block_U1084 ( .A(aes_core_round_key[48]), .B(
        aes_core_enc_block_n1426), .Y(aes_core_enc_block_n832) );
  AOI222X1 aes_core_enc_block_U1083 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[16]), .B0(aes_core_enc_block_n51), .B1(
        aes_core_enc_block_n832), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n833), .Y(aes_core_enc_block_n831) );
  XNOR2X1 aes_core_enc_block_U1082 ( .A(aes_core_round_key[48]), .B(Din[48]), 
        .Y(aes_core_enc_block_n830) );
  OAI221X1 aes_core_enc_block_U1081 ( .A0(aes_core_enc_block_n830), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1427), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n831), .Y(
        aes_core_enc_block_n1289) );
  XNOR2X1 aes_core_enc_block_U1080 ( .A(aes_core_round_key[16]), .B(
        aes_core_enc_block_n1424), .Y(aes_core_enc_block_n1071) );
  AOI222X1 aes_core_enc_block_U1079 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[16]), .B0(aes_core_enc_block_n58), .B1(
        aes_core_enc_block_n1071), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n1072), .Y(aes_core_enc_block_n1070) );
  XNOR2X1 aes_core_enc_block_U1078 ( .A(aes_core_round_key[16]), .B(Din[16]), 
        .Y(aes_core_enc_block_n1069) );
  OAI221X1 aes_core_enc_block_U1077 ( .A0(aes_core_enc_block_n1069), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1426), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1070), .Y(
        aes_core_enc_block_n1321) );
  XOR2X1 aes_core_enc_block_U1076 ( .A(aes_core_enc_block_n977), .B(
        aes_core_enc_block_n978), .Y(aes_core_enc_block_n974) );
  OAI2BB2X1 aes_core_enc_block_U1075 ( .B0(aes_core_enc_block_n1389), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n115), .A1N(Din[28]), 
        .Y(aes_core_enc_block_n975) );
  AOI222X1 aes_core_enc_block_U1074 ( .A0(aes_core_enc_block_n119), .A1(
        aes_core_enc_block_n974), .B0(aes_core_enc_block_n975), .B1(
        aes_core_enc_block_n167), .C0(aes_core_round_key[28]), .C1(
        aes_core_enc_block_n976), .Y(aes_core_enc_block_n973) );
  OAI221X1 aes_core_enc_block_U1073 ( .A0(aes_core_enc_block_n158), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1389), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n973), .Y(
        aes_core_enc_block_n1309) );
  XOR2X1 aes_core_enc_block_U1072 ( .A(aes_core_enc_block_n1004), .B(
        aes_core_enc_block_n1005), .Y(aes_core_enc_block_n1001) );
  OAI2BB2X1 aes_core_enc_block_U1071 ( .B0(aes_core_enc_block_n1438), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n116), .A1N(Din[25]), 
        .Y(aes_core_enc_block_n1002) );
  AOI222X1 aes_core_enc_block_U1070 ( .A0(aes_core_enc_block_n119), .A1(
        aes_core_enc_block_n1001), .B0(aes_core_enc_block_n1002), .B1(
        aes_core_enc_block_n170), .C0(aes_core_round_key[25]), .C1(
        aes_core_enc_block_n1003), .Y(aes_core_enc_block_n1000) );
  OAI221X1 aes_core_enc_block_U1069 ( .A0(aes_core_enc_block_n163), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1438), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1000), .Y(
        aes_core_enc_block_n1312) );
  OAI2BB2X1 aes_core_enc_block_U1068 ( .B0(aes_core_enc_block_n1447), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n116), .A1N(Din[26]), 
        .Y(aes_core_enc_block_n994) );
  XOR2X1 aes_core_enc_block_U1067 ( .A(aes_core_enc_block_n996), .B(
        aes_core_enc_block_n997), .Y(aes_core_enc_block_n993) );
  AOI222X1 aes_core_enc_block_U1066 ( .A0(aes_core_enc_block_n118), .A1(
        aes_core_enc_block_n993), .B0(aes_core_enc_block_n994), .B1(
        aes_core_enc_block_n169), .C0(aes_core_round_key[26]), .C1(
        aes_core_enc_block_n995), .Y(aes_core_enc_block_n992) );
  OAI221X1 aes_core_enc_block_U1065 ( .A0(aes_core_enc_block_n161), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1447), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n992), .Y(
        aes_core_enc_block_n1311) );
  XNOR2X1 aes_core_enc_block_U1064 ( .A(aes_core_round_key[107]), .B(
        aes_core_enc_block_n1348), .Y(aes_core_enc_block_n391) );
  AOI222X1 aes_core_enc_block_U1063 ( .A0(aes_core_new_sboxw[11]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n34), .B1(
        aes_core_enc_block_n391), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n392), .Y(aes_core_enc_block_n390) );
  XNOR2X1 aes_core_enc_block_U1062 ( .A(aes_core_round_key[107]), .B(Din[107]), 
        .Y(aes_core_enc_block_n389) );
  OAI221X1 aes_core_enc_block_U1061 ( .A0(aes_core_enc_block_n389), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n190), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n390), .Y(
        aes_core_enc_block_n1231) );
  XNOR2X1 aes_core_enc_block_U1060 ( .A(aes_core_round_key[40]), .B(
        aes_core_enc_block_n1422), .Y(aes_core_enc_block_n884) );
  AOI222X1 aes_core_enc_block_U1059 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[8]), .B0(aes_core_enc_block_n55), .B1(
        aes_core_enc_block_n884), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n885), .Y(aes_core_enc_block_n883) );
  XNOR2X1 aes_core_enc_block_U1058 ( .A(aes_core_round_key[40]), .B(Din[40]), 
        .Y(aes_core_enc_block_n882) );
  OAI221X1 aes_core_enc_block_U1057 ( .A0(aes_core_enc_block_n882), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1423), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n883), .Y(
        aes_core_enc_block_n1297) );
  XNOR2X1 aes_core_enc_block_U1056 ( .A(aes_core_round_key[112]), .B(
        aes_core_enc_block_n1430), .Y(aes_core_enc_block_n359) );
  AOI222X1 aes_core_enc_block_U1055 ( .A0(aes_core_new_sboxw[16]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n30), .B1(
        aes_core_enc_block_n359), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n360), .Y(aes_core_enc_block_n358) );
  XNOR2X1 aes_core_enc_block_U1054 ( .A(aes_core_round_key[112]), .B(Din[112]), 
        .Y(aes_core_enc_block_n357) );
  OAI221X1 aes_core_enc_block_U1053 ( .A0(aes_core_enc_block_n357), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1424), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n358), .Y(
        aes_core_enc_block_n1226) );
  XNOR2X1 aes_core_enc_block_U1052 ( .A(aes_core_round_key[114]), .B(
        aes_core_enc_block_n1444), .Y(aes_core_enc_block_n344) );
  AOI222X1 aes_core_enc_block_U1051 ( .A0(aes_core_new_sboxw[18]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n31), .B1(
        aes_core_enc_block_n344), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n345), .Y(aes_core_enc_block_n343) );
  XNOR2X1 aes_core_enc_block_U1050 ( .A(aes_core_round_key[114]), .B(Din[114]), 
        .Y(aes_core_enc_block_n342) );
  OAI221X1 aes_core_enc_block_U1049 ( .A0(aes_core_enc_block_n342), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1446), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n343), .Y(
        aes_core_enc_block_n1224) );
  XOR2X1 aes_core_enc_block_U1048 ( .A(aes_core_enc_block_n275), .B(
        aes_core_enc_block_n276), .Y(aes_core_enc_block_n272) );
  OAI2BB2X1 aes_core_enc_block_U1047 ( .B0(aes_core_enc_block_n1449), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n110), .A1N(Din[123]), 
        .Y(aes_core_enc_block_n273) );
  AOI222X1 aes_core_enc_block_U1046 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n272), .B0(aes_core_enc_block_n273), .B1(
        aes_core_enc_block_n136), .C0(aes_core_round_key[123]), .C1(
        aes_core_enc_block_n274), .Y(aes_core_enc_block_n271) );
  OAI221X1 aes_core_enc_block_U1045 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n162), .B0(aes_core_enc_block_n1449), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n271), .Y(
        aes_core_enc_block_n1215) );
  OAI2BB2X1 aes_core_enc_block_U1044 ( .B0(aes_core_enc_block_n1395), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n113), .A1N(Din[56]), 
        .Y(aes_core_enc_block_n772) );
  XOR2X1 aes_core_enc_block_U1043 ( .A(aes_core_enc_block_n774), .B(
        aes_core_enc_block_n775), .Y(aes_core_enc_block_n771) );
  AOI222X1 aes_core_enc_block_U1042 ( .A0(aes_core_enc_block_n119), .A1(
        aes_core_enc_block_n771), .B0(aes_core_enc_block_n772), .B1(
        aes_core_enc_block_n155), .C0(aes_core_round_key[56]), .C1(
        aes_core_enc_block_n773), .Y(aes_core_enc_block_n770) );
  OAI221X1 aes_core_enc_block_U1041 ( .A0(aes_core_enc_block_n164), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1395), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n770), .Y(
        aes_core_enc_block_n1281) );
  OAI2BB2X1 aes_core_enc_block_U1040 ( .B0(aes_core_enc_block_n1441), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n114), .A1N(Din[58]), 
        .Y(aes_core_enc_block_n755) );
  XOR2X1 aes_core_enc_block_U1039 ( .A(aes_core_enc_block_n757), .B(
        aes_core_enc_block_n758), .Y(aes_core_enc_block_n754) );
  AOI222X1 aes_core_enc_block_U1038 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n754), .B0(aes_core_enc_block_n755), .B1(
        aes_core_enc_block_n153), .C0(aes_core_round_key[58]), .C1(
        aes_core_enc_block_n756), .Y(aes_core_enc_block_n753) );
  OAI221X1 aes_core_enc_block_U1037 ( .A0(aes_core_enc_block_n161), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1441), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n753), .Y(
        aes_core_enc_block_n1279) );
  XOR2X1 aes_core_enc_block_U1036 ( .A(aes_core_enc_block_n748), .B(
        aes_core_enc_block_n749), .Y(aes_core_enc_block_n745) );
  OAI2BB2X1 aes_core_enc_block_U1035 ( .B0(aes_core_enc_block_n1453), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n113), .A1N(Din[59]), 
        .Y(aes_core_enc_block_n746) );
  AOI222X1 aes_core_enc_block_U1034 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n745), .B0(aes_core_enc_block_n746), .B1(
        aes_core_enc_block_n152), .C0(aes_core_round_key[59]), .C1(
        aes_core_enc_block_n747), .Y(aes_core_enc_block_n744) );
  OAI221X1 aes_core_enc_block_U1033 ( .A0(aes_core_enc_block_n162), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1453), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n744), .Y(
        aes_core_enc_block_n1278) );
  OAI2BB2X1 aes_core_enc_block_U1032 ( .B0(aes_core_enc_block_n1425), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n107), .A1N(Din[24]), 
        .Y(aes_core_enc_block_n1011) );
  XOR2X1 aes_core_enc_block_U1031 ( .A(aes_core_enc_block_n1013), .B(
        aes_core_enc_block_n1014), .Y(aes_core_enc_block_n1010) );
  AOI222X1 aes_core_enc_block_U1030 ( .A0(aes_core_enc_block_n120), .A1(
        aes_core_enc_block_n1010), .B0(aes_core_enc_block_n1011), .B1(
        aes_core_enc_block_n171), .C0(aes_core_round_key[24]), .C1(
        aes_core_enc_block_n1012), .Y(aes_core_enc_block_n1009) );
  OAI221X1 aes_core_enc_block_U1029 ( .A0(aes_core_enc_block_n164), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1425), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1009), .Y(
        aes_core_enc_block_n1313) );
  XNOR2X1 aes_core_enc_block_U1028 ( .A(aes_core_round_key[53]), .B(
        aes_core_enc_block_n1405), .Y(aes_core_enc_block_n794) );
  AOI222X1 aes_core_enc_block_U1027 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[21]), .B0(aes_core_enc_block_n49), .B1(
        aes_core_enc_block_n794), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n795), .Y(aes_core_enc_block_n793) );
  XNOR2X1 aes_core_enc_block_U1026 ( .A(aes_core_round_key[53]), .B(Din[53]), 
        .Y(aes_core_enc_block_n792) );
  OAI221X1 aes_core_enc_block_U1025 ( .A0(aes_core_enc_block_n792), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1406), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n793), .Y(
        aes_core_enc_block_n1284) );
  XNOR2X1 aes_core_enc_block_U1024 ( .A(aes_core_round_key[49]), .B(
        aes_core_enc_block_n1439), .Y(aes_core_enc_block_n824) );
  AOI222X1 aes_core_enc_block_U1023 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[17]), .B0(aes_core_enc_block_n50), .B1(
        aes_core_enc_block_n824), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n825), .Y(aes_core_enc_block_n823) );
  XNOR2X1 aes_core_enc_block_U1022 ( .A(aes_core_round_key[49]), .B(Din[49]), 
        .Y(aes_core_enc_block_n822) );
  OAI221X1 aes_core_enc_block_U1021 ( .A0(aes_core_enc_block_n822), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1431), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n823), .Y(
        aes_core_enc_block_n1288) );
  XNOR2X1 aes_core_enc_block_U1020 ( .A(aes_core_round_key[21]), .B(
        aes_core_enc_block_n1378), .Y(aes_core_enc_block_n1033) );
  AOI222X1 aes_core_enc_block_U1019 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[21]), .B0(aes_core_enc_block_n58), .B1(
        aes_core_enc_block_n1033), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n1034), .Y(aes_core_enc_block_n1032) );
  XNOR2X1 aes_core_enc_block_U1018 ( .A(aes_core_round_key[21]), .B(Din[21]), 
        .Y(aes_core_enc_block_n1031) );
  OAI221X1 aes_core_enc_block_U1017 ( .A0(aes_core_enc_block_n1031), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1405), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1032), .Y(
        aes_core_enc_block_n1316) );
  XNOR2X1 aes_core_enc_block_U1016 ( .A(aes_core_round_key[17]), .B(
        aes_core_enc_block_n1435), .Y(aes_core_enc_block_n1063) );
  AOI222X1 aes_core_enc_block_U1015 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[17]), .B0(aes_core_enc_block_n59), .B1(
        aes_core_enc_block_n1063), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n1064), .Y(aes_core_enc_block_n1062) );
  XNOR2X1 aes_core_enc_block_U1014 ( .A(aes_core_round_key[17]), .B(Din[17]), 
        .Y(aes_core_enc_block_n1061) );
  OAI221X1 aes_core_enc_block_U1013 ( .A0(aes_core_enc_block_n1061), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1439), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1062), .Y(
        aes_core_enc_block_n1320) );
  XOR2X1 aes_core_enc_block_U1012 ( .A(aes_core_enc_block_n524), .B(
        aes_core_enc_block_n525), .Y(aes_core_enc_block_n521) );
  OAI2BB2X1 aes_core_enc_block_U1011 ( .B0(aes_core_enc_block_n1432), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n112), .A1N(Din[89]), 
        .Y(aes_core_enc_block_n522) );
  AOI222X1 aes_core_enc_block_U1010 ( .A0(aes_core_enc_block_n120), .A1(
        aes_core_enc_block_n521), .B0(aes_core_enc_block_n522), .B1(
        aes_core_enc_block_n146), .C0(aes_core_round_key[89]), .C1(
        aes_core_enc_block_n523), .Y(aes_core_enc_block_n520) );
  OAI221X1 aes_core_enc_block_U1009 ( .A0(aes_core_enc_block_n163), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1432), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n520), .Y(
        aes_core_enc_block_n1248) );
  OAI2BB2X1 aes_core_enc_block_U1008 ( .B0(aes_core_enc_block_n1443), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n108), .A1N(Din[90]), 
        .Y(aes_core_enc_block_n514) );
  XOR2X1 aes_core_enc_block_U1007 ( .A(aes_core_enc_block_n516), .B(
        aes_core_enc_block_n517), .Y(aes_core_enc_block_n513) );
  AOI222X1 aes_core_enc_block_U1006 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n513), .B0(aes_core_enc_block_n514), .B1(
        aes_core_enc_block_n145), .C0(aes_core_round_key[90]), .C1(
        aes_core_enc_block_n515), .Y(aes_core_enc_block_n512) );
  OAI221X1 aes_core_enc_block_U1005 ( .A0(aes_core_enc_block_n161), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1443), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n512), .Y(
        aes_core_enc_block_n1247) );
  XNOR2X1 aes_core_enc_block_U1004 ( .A(aes_core_round_key[96]), .B(
        aes_core_enc_block_n947), .Y(aes_core_enc_block_n1188) );
  AOI222X1 aes_core_enc_block_U1003 ( .A0(aes_core_new_sboxw[0]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n65), .B1(
        aes_core_enc_block_n1188), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n1189), .Y(aes_core_enc_block_n1187) );
  XNOR2X1 aes_core_enc_block_U1002 ( .A(aes_core_round_key[96]), .B(Din[96]), 
        .Y(aes_core_enc_block_n1186) );
  OAI221X1 aes_core_enc_block_U1001 ( .A0(aes_core_enc_block_n1186), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n187), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n1187), .Y(
        aes_core_enc_block_n1338) );
  XNOR2X1 aes_core_enc_block_U1000 ( .A(aes_core_round_key[32]), .B(
        aes_core_enc_block_n1362), .Y(aes_core_enc_block_n942) );
  AOI222X1 aes_core_enc_block_U999 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[0]), .B0(aes_core_enc_block_n56), .B1(
        aes_core_enc_block_n942), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n943), .Y(aes_core_enc_block_n941) );
  XNOR2X1 aes_core_enc_block_U998 ( .A(aes_core_round_key[32]), .B(Din[32]), 
        .Y(aes_core_enc_block_n940) );
  OAI221X1 aes_core_enc_block_U997 ( .A0(aes_core_enc_block_n940), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1396), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n941), .Y(
        aes_core_enc_block_n1305) );
  XNOR2X1 aes_core_enc_block_U996 ( .A(aes_core_round_key[0]), .B(
        aes_core_enc_block_n1396), .Y(aes_core_enc_block_n1181) );
  AOI222X1 aes_core_enc_block_U995 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[0]), .B0(aes_core_enc_block_n53), .B1(
        aes_core_enc_block_n1181), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1182), .Y(aes_core_enc_block_n1180) );
  XNOR2X1 aes_core_enc_block_U994 ( .A(aes_core_round_key[0]), .B(Din[0]), .Y(
        aes_core_enc_block_n1179) );
  OAI221X1 aes_core_enc_block_U993 ( .A0(aes_core_enc_block_n1179), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n947), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1180), .Y(
        aes_core_enc_block_n1337) );
  OAI2BB2X1 aes_core_enc_block_U992 ( .B0(aes_core_enc_block_n1379), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n115), .A1N(Din[29]), 
        .Y(aes_core_enc_block_n967) );
  XOR2X1 aes_core_enc_block_U991 ( .A(aes_core_enc_block_n969), .B(
        aes_core_enc_block_n970), .Y(aes_core_enc_block_n966) );
  AOI222X1 aes_core_enc_block_U990 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n966), .B0(aes_core_enc_block_n967), .B1(
        aes_core_enc_block_n166), .C0(aes_core_round_key[29]), .C1(
        aes_core_enc_block_n968), .Y(aes_core_enc_block_n965) );
  OAI221X1 aes_core_enc_block_U989 ( .A0(aes_core_enc_block_n160), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1379), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n965), .Y(
        aes_core_enc_block_n1308) );
  OAI2BB2X1 aes_core_enc_block_U988 ( .B0(aes_core_enc_block_n1380), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n115), .A1N(Din[30]), 
        .Y(aes_core_enc_block_n959) );
  XOR2X1 aes_core_enc_block_U987 ( .A(aes_core_enc_block_n961), .B(
        aes_core_enc_block_n962), .Y(aes_core_enc_block_n958) );
  AOI222X1 aes_core_enc_block_U986 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n958), .B0(aes_core_enc_block_n959), .B1(
        aes_core_enc_block_n165), .C0(aes_core_round_key[30]), .C1(
        aes_core_enc_block_n960), .Y(aes_core_enc_block_n957) );
  OAI221X1 aes_core_enc_block_U985 ( .A0(aes_core_enc_block_n157), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1380), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n957), .Y(
        aes_core_enc_block_n1307) );
  XNOR2X1 aes_core_enc_block_U984 ( .A(aes_core_round_key[85]), .B(
        aes_core_enc_block_n1406), .Y(aes_core_enc_block_n553) );
  AOI222X1 aes_core_enc_block_U983 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[21]), .B0(aes_core_enc_block_n39), .B1(
        aes_core_enc_block_n553), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n554), .Y(aes_core_enc_block_n552) );
  XNOR2X1 aes_core_enc_block_U982 ( .A(aes_core_round_key[85]), .B(Din[85]), 
        .Y(aes_core_enc_block_n551) );
  OAI221X1 aes_core_enc_block_U981 ( .A0(aes_core_enc_block_n551), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1407), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n552), .Y(
        aes_core_enc_block_n1252) );
  XNOR2X1 aes_core_enc_block_U980 ( .A(aes_core_round_key[80]), .B(
        aes_core_enc_block_n1427), .Y(aes_core_enc_block_n591) );
  AOI222X1 aes_core_enc_block_U979 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[16]), .B0(aes_core_enc_block_n40), .B1(
        aes_core_enc_block_n591), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n592), .Y(aes_core_enc_block_n590) );
  XNOR2X1 aes_core_enc_block_U978 ( .A(aes_core_round_key[80]), .B(Din[80]), 
        .Y(aes_core_enc_block_n589) );
  OAI221X1 aes_core_enc_block_U977 ( .A0(aes_core_enc_block_n589), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1430), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n590), .Y(
        aes_core_enc_block_n1257) );
  XNOR2X1 aes_core_enc_block_U976 ( .A(aes_core_round_key[81]), .B(
        aes_core_enc_block_n1431), .Y(aes_core_enc_block_n583) );
  AOI222X1 aes_core_enc_block_U975 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[17]), .B0(aes_core_enc_block_n41), .B1(
        aes_core_enc_block_n583), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n584), .Y(aes_core_enc_block_n582) );
  XNOR2X1 aes_core_enc_block_U974 ( .A(aes_core_round_key[81]), .B(Din[81]), 
        .Y(aes_core_enc_block_n581) );
  OAI221X1 aes_core_enc_block_U973 ( .A0(aes_core_enc_block_n581), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1433), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n582), .Y(
        aes_core_enc_block_n1256) );
  OAI2BB2X1 aes_core_enc_block_U972 ( .B0(aes_core_enc_block_n1429), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n107), .A1N(Din[88]), 
        .Y(aes_core_enc_block_n531) );
  XOR2X1 aes_core_enc_block_U971 ( .A(aes_core_enc_block_n533), .B(
        aes_core_enc_block_n534), .Y(aes_core_enc_block_n530) );
  AOI222X1 aes_core_enc_block_U970 ( .A0(aes_core_enc_block_n118), .A1(
        aes_core_enc_block_n530), .B0(aes_core_enc_block_n531), .B1(
        aes_core_enc_block_n147), .C0(aes_core_round_key[88]), .C1(
        aes_core_enc_block_n532), .Y(aes_core_enc_block_n529) );
  OAI221X1 aes_core_enc_block_U969 ( .A0(aes_core_enc_block_n164), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1429), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n529), .Y(
        aes_core_enc_block_n1249) );
  XOR2X1 aes_core_enc_block_U968 ( .A(aes_core_enc_block_n507), .B(
        aes_core_enc_block_n508), .Y(aes_core_enc_block_n504) );
  OAI2BB2X1 aes_core_enc_block_U967 ( .B0(aes_core_enc_block_n1452), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n111), .A1N(Din[91]), 
        .Y(aes_core_enc_block_n505) );
  AOI222X1 aes_core_enc_block_U966 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n504), .B0(aes_core_enc_block_n505), .B1(
        aes_core_enc_block_n144), .C0(aes_core_round_key[91]), .C1(
        aes_core_enc_block_n506), .Y(aes_core_enc_block_n503) );
  OAI221X1 aes_core_enc_block_U965 ( .A0(aes_core_enc_block_n162), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1452), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n503), .Y(
        aes_core_enc_block_n1246) );
  XOR2X1 aes_core_enc_block_U964 ( .A(aes_core_enc_block_n738), .B(
        aes_core_enc_block_n739), .Y(aes_core_enc_block_n735) );
  OAI2BB2X1 aes_core_enc_block_U963 ( .B0(aes_core_enc_block_n1391), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n113), .A1N(Din[60]), 
        .Y(aes_core_enc_block_n736) );
  AOI222X1 aes_core_enc_block_U962 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n735), .B0(aes_core_enc_block_n736), .B1(
        aes_core_enc_block_n151), .C0(aes_core_round_key[60]), .C1(
        aes_core_enc_block_n737), .Y(aes_core_enc_block_n734) );
  OAI221X1 aes_core_enc_block_U961 ( .A0(aes_core_enc_block_n158), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1391), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n734), .Y(
        aes_core_enc_block_n1277) );
  OAI2BB2X1 aes_core_enc_block_U960 ( .B0(aes_core_enc_block_n1392), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n110), .A1N(Din[61]), 
        .Y(aes_core_enc_block_n728) );
  XOR2X1 aes_core_enc_block_U959 ( .A(aes_core_enc_block_n730), .B(
        aes_core_enc_block_n731), .Y(aes_core_enc_block_n727) );
  AOI222X1 aes_core_enc_block_U958 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n727), .B0(aes_core_enc_block_n728), .B1(
        aes_core_enc_block_n150), .C0(aes_core_round_key[61]), .C1(
        aes_core_enc_block_n729), .Y(aes_core_enc_block_n726) );
  OAI221X1 aes_core_enc_block_U957 ( .A0(aes_core_enc_block_n160), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1392), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n726), .Y(
        aes_core_enc_block_n1276) );
  OAI2BB2X1 aes_core_enc_block_U956 ( .B0(aes_core_enc_block_n1393), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n112), .A1N(Din[62]), 
        .Y(aes_core_enc_block_n720) );
  XOR2X1 aes_core_enc_block_U955 ( .A(aes_core_enc_block_n722), .B(
        aes_core_enc_block_n723), .Y(aes_core_enc_block_n719) );
  AOI222X1 aes_core_enc_block_U954 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n719), .B0(aes_core_enc_block_n720), .B1(
        aes_core_enc_block_n149), .C0(aes_core_round_key[62]), .C1(
        aes_core_enc_block_n721), .Y(aes_core_enc_block_n718) );
  OAI221X1 aes_core_enc_block_U953 ( .A0(aes_core_enc_block_n157), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1393), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n718), .Y(
        aes_core_enc_block_n1275) );
  XOR2X1 aes_core_enc_block_U952 ( .A(aes_core_enc_block_n765), .B(
        aes_core_enc_block_n766), .Y(aes_core_enc_block_n762) );
  OAI2BB2X1 aes_core_enc_block_U951 ( .B0(aes_core_enc_block_n1440), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n114), .A1N(Din[57]), 
        .Y(aes_core_enc_block_n763) );
  AOI222X1 aes_core_enc_block_U950 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n762), .B0(aes_core_enc_block_n763), .B1(
        aes_core_enc_block_n154), .C0(aes_core_round_key[57]), .C1(
        aes_core_enc_block_n764), .Y(aes_core_enc_block_n761) );
  OAI221X1 aes_core_enc_block_U949 ( .A0(aes_core_enc_block_n163), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1440), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n761), .Y(
        aes_core_enc_block_n1280) );
  XNOR2X1 aes_core_enc_block_U948 ( .A(aes_core_round_key[108]), .B(
        aes_core_enc_block_n1377), .Y(aes_core_enc_block_n383) );
  AOI222X1 aes_core_enc_block_U947 ( .A0(aes_core_new_sboxw[12]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n33), .B1(
        aes_core_enc_block_n383), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n384), .Y(aes_core_enc_block_n382) );
  XNOR2X1 aes_core_enc_block_U946 ( .A(aes_core_round_key[108]), .B(Din[108]), 
        .Y(aes_core_enc_block_n381) );
  OAI221X1 aes_core_enc_block_U945 ( .A0(aes_core_enc_block_n381), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1349), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n382), .Y(
        aes_core_enc_block_n1230) );
  XNOR2X1 aes_core_enc_block_U944 ( .A(aes_core_round_key[106]), .B(
        aes_core_enc_block_n189), .Y(aes_core_enc_block_n398) );
  AOI222X1 aes_core_enc_block_U943 ( .A0(aes_core_new_sboxw[10]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n34), .B1(
        aes_core_enc_block_n398), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n399), .Y(aes_core_enc_block_n397) );
  XNOR2X1 aes_core_enc_block_U942 ( .A(aes_core_round_key[106]), .B(Din[106]), 
        .Y(aes_core_enc_block_n396) );
  OAI221X1 aes_core_enc_block_U941 ( .A0(aes_core_enc_block_n396), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1364), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n397), .Y(
        aes_core_enc_block_n1232) );
  XNOR2X1 aes_core_enc_block_U940 ( .A(aes_core_round_key[105]), .B(
        aes_core_enc_block_n1363), .Y(aes_core_enc_block_n404) );
  AOI222X1 aes_core_enc_block_U939 ( .A0(aes_core_new_sboxw[9]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n35), .B1(
        aes_core_enc_block_n404), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n405), .Y(aes_core_enc_block_n403) );
  XNOR2X1 aes_core_enc_block_U938 ( .A(aes_core_round_key[105]), .B(Din[105]), 
        .Y(aes_core_enc_block_n402) );
  OAI221X1 aes_core_enc_block_U937 ( .A0(aes_core_enc_block_n402), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1436), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n403), .Y(
        aes_core_enc_block_n1233) );
  XNOR2X1 aes_core_enc_block_U936 ( .A(aes_core_round_key[117]), .B(
        aes_core_enc_block_n1407), .Y(aes_core_enc_block_n321) );
  AOI222X1 aes_core_enc_block_U935 ( .A0(aes_core_new_sboxw[21]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n30), .B1(
        aes_core_enc_block_n321), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n322), .Y(aes_core_enc_block_n320) );
  XNOR2X1 aes_core_enc_block_U934 ( .A(aes_core_round_key[117]), .B(Din[117]), 
        .Y(aes_core_enc_block_n319) );
  OAI221X1 aes_core_enc_block_U933 ( .A0(aes_core_enc_block_n319), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1378), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n320), .Y(
        aes_core_enc_block_n1221) );
  XNOR2X1 aes_core_enc_block_U932 ( .A(aes_core_round_key[116]), .B(
        aes_core_enc_block_n1366), .Y(aes_core_enc_block_n328) );
  AOI222X1 aes_core_enc_block_U931 ( .A0(aes_core_new_sboxw[20]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n31), .B1(
        aes_core_enc_block_n328), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n329), .Y(aes_core_enc_block_n327) );
  XNOR2X1 aes_core_enc_block_U930 ( .A(aes_core_round_key[116]), .B(Din[116]), 
        .Y(aes_core_enc_block_n326) );
  OAI221X1 aes_core_enc_block_U929 ( .A0(aes_core_enc_block_n326), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1388), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n327), .Y(
        aes_core_enc_block_n1222) );
  XNOR2X1 aes_core_enc_block_U928 ( .A(aes_core_round_key[118]), .B(
        aes_core_enc_block_n1414), .Y(aes_core_enc_block_n314) );
  AOI222X1 aes_core_enc_block_U927 ( .A0(aes_core_new_sboxw[22]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n29), .B1(
        aes_core_enc_block_n314), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n315), .Y(aes_core_enc_block_n313) );
  XNOR2X1 aes_core_enc_block_U926 ( .A(aes_core_round_key[118]), .B(Din[118]), 
        .Y(aes_core_enc_block_n312) );
  OAI221X1 aes_core_enc_block_U925 ( .A0(aes_core_enc_block_n312), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1410), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n313), .Y(
        aes_core_enc_block_n1220) );
  XNOR2X1 aes_core_enc_block_U924 ( .A(aes_core_round_key[113]), .B(
        aes_core_enc_block_n1433), .Y(aes_core_enc_block_n351) );
  AOI222X1 aes_core_enc_block_U923 ( .A0(aes_core_new_sboxw[17]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n31), .B1(
        aes_core_enc_block_n351), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n352), .Y(aes_core_enc_block_n350) );
  XNOR2X1 aes_core_enc_block_U922 ( .A(aes_core_round_key[113]), .B(Din[113]), 
        .Y(aes_core_enc_block_n349) );
  OAI221X1 aes_core_enc_block_U921 ( .A0(aes_core_enc_block_n349), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1435), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n350), .Y(
        aes_core_enc_block_n1225) );
  XOR2X1 aes_core_enc_block_U920 ( .A(aes_core_enc_block_n265), .B(
        aes_core_enc_block_n266), .Y(aes_core_enc_block_n262) );
  OAI2BB2X1 aes_core_enc_block_U919 ( .B0(aes_core_enc_block_n1387), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n110), .A1N(Din[124]), 
        .Y(aes_core_enc_block_n263) );
  AOI222X1 aes_core_enc_block_U918 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n262), .B0(aes_core_enc_block_n263), .B1(
        aes_core_enc_block_n135), .C0(aes_core_round_key[124]), .C1(
        aes_core_enc_block_n264), .Y(aes_core_enc_block_n261) );
  OAI221X1 aes_core_enc_block_U917 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n158), .B0(aes_core_enc_block_n1387), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n261), .Y(
        aes_core_enc_block_n1214) );
  XOR2X1 aes_core_enc_block_U916 ( .A(aes_core_enc_block_n292), .B(
        aes_core_enc_block_n293), .Y(aes_core_enc_block_n289) );
  OAI2BB2X1 aes_core_enc_block_U915 ( .B0(aes_core_enc_block_n1434), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n108), .A1N(Din[121]), 
        .Y(aes_core_enc_block_n290) );
  AOI222X1 aes_core_enc_block_U914 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n289), .B0(aes_core_enc_block_n290), .B1(
        aes_core_enc_block_n138), .C0(aes_core_round_key[121]), .C1(
        aes_core_enc_block_n291), .Y(aes_core_enc_block_n288) );
  OAI221X1 aes_core_enc_block_U913 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n163), .B0(aes_core_enc_block_n1434), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n288), .Y(
        aes_core_enc_block_n1217) );
  OAI2BB2X1 aes_core_enc_block_U912 ( .B0(aes_core_enc_block_n1445), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n107), .A1N(Din[122]), 
        .Y(aes_core_enc_block_n282) );
  XOR2X1 aes_core_enc_block_U911 ( .A(aes_core_enc_block_n284), .B(
        aes_core_enc_block_n285), .Y(aes_core_enc_block_n281) );
  AOI222X1 aes_core_enc_block_U910 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n281), .B0(aes_core_enc_block_n282), .B1(
        aes_core_enc_block_n137), .C0(aes_core_round_key[122]), .C1(
        aes_core_enc_block_n283), .Y(aes_core_enc_block_n280) );
  OAI221X1 aes_core_enc_block_U909 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n161), .B0(aes_core_enc_block_n1445), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n280), .Y(
        aes_core_enc_block_n1216) );
  XNOR2X1 aes_core_enc_block_U908 ( .A(aes_core_round_key[104]), .B(
        aes_core_enc_block_n1423), .Y(aes_core_enc_block_n411) );
  AOI222X1 aes_core_enc_block_U907 ( .A0(aes_core_new_sboxw[8]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n35), .B1(
        aes_core_enc_block_n411), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n412), .Y(aes_core_enc_block_n410) );
  XNOR2X1 aes_core_enc_block_U906 ( .A(aes_core_round_key[104]), .B(Din[104]), 
        .Y(aes_core_enc_block_n409) );
  OAI221X1 aes_core_enc_block_U905 ( .A0(aes_core_enc_block_n409), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1422), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n410), .Y(
        aes_core_enc_block_n1234) );
  OAI2BB2X1 aes_core_enc_block_U904 ( .B0(aes_core_enc_block_n1421), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n107), .A1N(Din[120]), 
        .Y(aes_core_enc_block_n299) );
  XOR2X1 aes_core_enc_block_U903 ( .A(aes_core_enc_block_n301), .B(
        aes_core_enc_block_n302), .Y(aes_core_enc_block_n298) );
  AOI222X1 aes_core_enc_block_U902 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n298), .B0(aes_core_enc_block_n299), .B1(
        aes_core_enc_block_n139), .C0(aes_core_round_key[120]), .C1(
        aes_core_enc_block_n300), .Y(aes_core_enc_block_n297) );
  OAI221X1 aes_core_enc_block_U901 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n164), .B0(aes_core_enc_block_n1421), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n297), .Y(
        aes_core_enc_block_n1218) );
  OAI2BB2X1 aes_core_enc_block_U900 ( .B0(aes_core_enc_block_n1413), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n111), .A1N(Din[94]), 
        .Y(aes_core_enc_block_n479) );
  XOR2X1 aes_core_enc_block_U899 ( .A(aes_core_enc_block_n481), .B(
        aes_core_enc_block_n482), .Y(aes_core_enc_block_n478) );
  AOI222X1 aes_core_enc_block_U898 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n478), .B0(aes_core_enc_block_n479), .B1(
        aes_core_enc_block_n141), .C0(aes_core_round_key[94]), .C1(
        aes_core_enc_block_n480), .Y(aes_core_enc_block_n477) );
  OAI221X1 aes_core_enc_block_U897 ( .A0(aes_core_enc_block_n157), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1413), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n477), .Y(
        aes_core_enc_block_n1243) );
  XNOR2X1 aes_core_enc_block_U896 ( .A(aes_core_round_key[99]), .B(
        aes_core_enc_block_n1455), .Y(aes_core_enc_block_n446) );
  AOI222X1 aes_core_enc_block_U895 ( .A0(aes_core_new_sboxw[3]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n38), .B1(
        aes_core_enc_block_n446), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n447), .Y(aes_core_enc_block_n445) );
  XNOR2X1 aes_core_enc_block_U894 ( .A(aes_core_round_key[99]), .B(Din[99]), 
        .Y(aes_core_enc_block_n444) );
  OAI221X1 aes_core_enc_block_U893 ( .A0(aes_core_enc_block_n444), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1385), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n445), .Y(
        aes_core_enc_block_n1239) );
  XNOR2X1 aes_core_enc_block_U892 ( .A(aes_core_round_key[98]), .B(
        aes_core_enc_block_n1457), .Y(aes_core_enc_block_n454) );
  AOI222X1 aes_core_enc_block_U891 ( .A0(aes_core_new_sboxw[2]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n38), .B1(
        aes_core_enc_block_n454), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n455), .Y(aes_core_enc_block_n453) );
  XNOR2X1 aes_core_enc_block_U890 ( .A(aes_core_round_key[98]), .B(Din[98]), 
        .Y(aes_core_enc_block_n452) );
  OAI221X1 aes_core_enc_block_U889 ( .A0(aes_core_enc_block_n452), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1398), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n453), .Y(
        aes_core_enc_block_n1240) );
  XNOR2X1 aes_core_enc_block_U888 ( .A(aes_core_round_key[64]), .B(
        aes_core_enc_block_n187), .Y(aes_core_enc_block_n701) );
  AOI222X1 aes_core_enc_block_U887 ( .A0(aes_core_new_sboxw[0]), .A1(
        aes_core_enc_block_n9), .B0(aes_core_enc_block_n48), .B1(
        aes_core_enc_block_n701), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n702), .Y(aes_core_enc_block_n700) );
  XNOR2X1 aes_core_enc_block_U886 ( .A(aes_core_round_key[64]), .B(Din[64]), 
        .Y(aes_core_enc_block_n699) );
  OAI221X1 aes_core_enc_block_U885 ( .A0(aes_core_enc_block_n699), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1362), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n700), .Y(
        aes_core_enc_block_n1273) );
  XNOR2X1 aes_core_enc_block_U884 ( .A(aes_core_round_key[72]), .B(
        aes_core_enc_block_n1428), .Y(aes_core_enc_block_n643) );
  AOI222X1 aes_core_enc_block_U883 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[8]), .B0(aes_core_enc_block_n44), .B1(
        aes_core_enc_block_n643), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n644), .Y(aes_core_enc_block_n642) );
  XNOR2X1 aes_core_enc_block_U882 ( .A(aes_core_round_key[72]), .B(Din[72]), 
        .Y(aes_core_enc_block_n641) );
  OAI221X1 aes_core_enc_block_U881 ( .A0(aes_core_enc_block_n641), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1372), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n642), .Y(
        aes_core_enc_block_n1265) );
  XOR2X1 aes_core_enc_block_U880 ( .A(aes_core_enc_block_n497), .B(
        aes_core_enc_block_n498), .Y(aes_core_enc_block_n494) );
  OAI2BB2X1 aes_core_enc_block_U879 ( .B0(aes_core_enc_block_n1402), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n111), .A1N(Din[92]), 
        .Y(aes_core_enc_block_n495) );
  AOI222X1 aes_core_enc_block_U878 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n494), .B0(aes_core_enc_block_n495), .B1(
        aes_core_enc_block_n143), .C0(aes_core_round_key[92]), .C1(
        aes_core_enc_block_n496), .Y(aes_core_enc_block_n493) );
  OAI221X1 aes_core_enc_block_U877 ( .A0(aes_core_enc_block_n158), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1402), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n493), .Y(
        aes_core_enc_block_n1245) );
  OAI2BB2X1 aes_core_enc_block_U876 ( .B0(aes_core_enc_block_n1403), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n111), .A1N(Din[93]), 
        .Y(aes_core_enc_block_n487) );
  XOR2X1 aes_core_enc_block_U875 ( .A(aes_core_enc_block_n489), .B(
        aes_core_enc_block_n490), .Y(aes_core_enc_block_n486) );
  AOI222X1 aes_core_enc_block_U874 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n486), .B0(aes_core_enc_block_n487), .B1(
        aes_core_enc_block_n142), .C0(aes_core_round_key[93]), .C1(
        aes_core_enc_block_n488), .Y(aes_core_enc_block_n485) );
  OAI221X1 aes_core_enc_block_U873 ( .A0(aes_core_enc_block_n160), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1403), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n485), .Y(
        aes_core_enc_block_n1244) );
  OAI2BB2X1 aes_core_enc_block_U872 ( .B0(aes_core_enc_block_n1408), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n110), .A1N(Din[125]), 
        .Y(aes_core_enc_block_n255) );
  XOR2X1 aes_core_enc_block_U871 ( .A(aes_core_enc_block_n257), .B(
        aes_core_enc_block_n258), .Y(aes_core_enc_block_n254) );
  AOI222X1 aes_core_enc_block_U870 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n254), .B0(aes_core_enc_block_n255), .B1(
        aes_core_enc_block_n134), .C0(aes_core_round_key[125]), .C1(
        aes_core_enc_block_n256), .Y(aes_core_enc_block_n253) );
  OAI221X1 aes_core_enc_block_U869 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n160), .B0(aes_core_enc_block_n1408), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n253), .Y(
        aes_core_enc_block_n1213) );
  OAI2BB2X1 aes_core_enc_block_U868 ( .B0(aes_core_enc_block_n1409), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n108), .A1N(Din[126]), 
        .Y(aes_core_enc_block_n247) );
  XOR2X1 aes_core_enc_block_U867 ( .A(aes_core_enc_block_n249), .B(
        aes_core_enc_block_n250), .Y(aes_core_enc_block_n246) );
  AOI222X1 aes_core_enc_block_U866 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n246), .B0(aes_core_enc_block_n247), .B1(
        aes_core_enc_block_n133), .C0(aes_core_round_key[126]), .C1(
        aes_core_enc_block_n248), .Y(aes_core_enc_block_n245) );
  OAI221X1 aes_core_enc_block_U865 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n157), .B0(aes_core_enc_block_n1409), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n245), .Y(
        aes_core_enc_block_n1212) );
  XNOR2X1 aes_core_enc_block_U864 ( .A(aes_core_round_key[8]), .B(
        aes_core_enc_block_n1372), .Y(aes_core_enc_block_n1123) );
  AOI222X1 aes_core_enc_block_U863 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[8]), .B0(aes_core_enc_block_n63), .B1(
        aes_core_enc_block_n1123), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1124), .Y(aes_core_enc_block_n1122) );
  XNOR2X1 aes_core_enc_block_U862 ( .A(aes_core_round_key[8]), .B(Din[8]), .Y(
        aes_core_enc_block_n1121) );
  OAI221X1 aes_core_enc_block_U861 ( .A0(aes_core_enc_block_n1121), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1428), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1122), .Y(
        aes_core_enc_block_n1329) );
  XNOR2X1 aes_core_enc_block_U860 ( .A(aes_core_round_key[110]), .B(
        aes_core_enc_block_n1356), .Y(aes_core_enc_block_n371) );
  AOI222X1 aes_core_enc_block_U859 ( .A0(aes_core_new_sboxw[14]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n32), .B1(
        aes_core_enc_block_n371), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n372), .Y(aes_core_enc_block_n370) );
  XNOR2X1 aes_core_enc_block_U858 ( .A(aes_core_round_key[110]), .B(Din[110]), 
        .Y(aes_core_enc_block_n369) );
  OAI221X1 aes_core_enc_block_U857 ( .A0(aes_core_enc_block_n369), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n196), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n370), .Y(
        aes_core_enc_block_n1228) );
  XNOR2X1 aes_core_enc_block_U856 ( .A(aes_core_round_key[101]), .B(
        aes_core_enc_block_n195), .Y(aes_core_enc_block_n431) );
  AOI222X1 aes_core_enc_block_U855 ( .A0(aes_core_new_sboxw[5]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n37), .B1(
        aes_core_enc_block_n431), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n432), .Y(aes_core_enc_block_n430) );
  XNOR2X1 aes_core_enc_block_U854 ( .A(aes_core_round_key[101]), .B(Din[101]), 
        .Y(aes_core_enc_block_n429) );
  OAI221X1 aes_core_enc_block_U853 ( .A0(aes_core_enc_block_n429), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1354), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n430), .Y(
        aes_core_enc_block_n1237) );
  XNOR2X1 aes_core_enc_block_U852 ( .A(aes_core_round_key[102]), .B(
        aes_core_enc_block_n240), .Y(aes_core_enc_block_n424) );
  AOI222X1 aes_core_enc_block_U851 ( .A0(aes_core_new_sboxw[6]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n36), .B1(
        aes_core_enc_block_n424), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n425), .Y(aes_core_enc_block_n423) );
  XNOR2X1 aes_core_enc_block_U850 ( .A(aes_core_round_key[102]), .B(Din[102]), 
        .Y(aes_core_enc_block_n422) );
  OAI221X1 aes_core_enc_block_U849 ( .A0(aes_core_enc_block_n422), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1357), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n423), .Y(
        aes_core_enc_block_n1236) );
  XNOR2X1 aes_core_enc_block_U848 ( .A(aes_core_round_key[100]), .B(
        aes_core_enc_block_n192), .Y(aes_core_enc_block_n438) );
  AOI222X1 aes_core_enc_block_U847 ( .A0(aes_core_new_sboxw[4]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n37), .B1(
        aes_core_enc_block_n438), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n439), .Y(aes_core_enc_block_n437) );
  XNOR2X1 aes_core_enc_block_U846 ( .A(aes_core_round_key[100]), .B(Din[100]), 
        .Y(aes_core_enc_block_n436) );
  OAI221X1 aes_core_enc_block_U845 ( .A0(aes_core_enc_block_n436), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1367), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n437), .Y(
        aes_core_enc_block_n1238) );
  XNOR2X1 aes_core_enc_block_U844 ( .A(aes_core_round_key[97]), .B(
        aes_core_enc_block_n1397), .Y(aes_core_enc_block_n461) );
  AOI222X1 aes_core_enc_block_U843 ( .A0(aes_core_new_sboxw[1]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n39), .B1(
        aes_core_enc_block_n461), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n462), .Y(aes_core_enc_block_n460) );
  XNOR2X1 aes_core_enc_block_U842 ( .A(aes_core_round_key[97]), .B(Din[97]), 
        .Y(aes_core_enc_block_n459) );
  OAI221X1 aes_core_enc_block_U841 ( .A0(aes_core_enc_block_n459), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1207), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n460), .Y(
        aes_core_enc_block_n1241) );
  XNOR2X1 aes_core_enc_block_U840 ( .A(aes_core_round_key[4]), .B(
        aes_core_enc_block_n1350), .Y(aes_core_enc_block_n1150) );
  AOI222X1 aes_core_enc_block_U839 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[4]), .B0(aes_core_enc_block_n63), .B1(
        aes_core_enc_block_n1150), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n1151), .Y(aes_core_enc_block_n1149) );
  XNOR2X1 aes_core_enc_block_U838 ( .A(aes_core_round_key[4]), .B(Din[4]), .Y(
        aes_core_enc_block_n1148) );
  OAI221X1 aes_core_enc_block_U837 ( .A0(aes_core_enc_block_n1148), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n192), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1149), .Y(
        aes_core_enc_block_n1333) );
  XNOR2X1 aes_core_enc_block_U836 ( .A(aes_core_round_key[38]), .B(
        aes_core_enc_block_n1358), .Y(aes_core_enc_block_n897) );
  AOI222X1 aes_core_enc_block_U835 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[6]), .B0(aes_core_enc_block_n54), .B1(
        aes_core_enc_block_n897), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n898), .Y(aes_core_enc_block_n896) );
  XNOR2X1 aes_core_enc_block_U834 ( .A(aes_core_round_key[38]), .B(Din[38]), 
        .Y(aes_core_enc_block_n895) );
  OAI221X1 aes_core_enc_block_U833 ( .A0(aes_core_enc_block_n895), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n232), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n896), .Y(
        aes_core_enc_block_n1299) );
  XNOR2X1 aes_core_enc_block_U832 ( .A(aes_core_round_key[6]), .B(
        aes_core_enc_block_n232), .Y(aes_core_enc_block_n1136) );
  AOI222X1 aes_core_enc_block_U831 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[6]), .B0(aes_core_enc_block_n62), .B1(
        aes_core_enc_block_n1136), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n1137), .Y(aes_core_enc_block_n1135) );
  XNOR2X1 aes_core_enc_block_U830 ( .A(aes_core_round_key[6]), .B(Din[6]), .Y(
        aes_core_enc_block_n1134) );
  OAI221X1 aes_core_enc_block_U829 ( .A0(aes_core_enc_block_n1134), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n240), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1135), .Y(
        aes_core_enc_block_n1331) );
  XNOR2X1 aes_core_enc_block_U828 ( .A(aes_core_round_key[36]), .B(
        aes_core_enc_block_n1352), .Y(aes_core_enc_block_n911) );
  AOI222X1 aes_core_enc_block_U827 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[4]), .B0(aes_core_enc_block_n55), .B1(
        aes_core_enc_block_n911), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n912), .Y(aes_core_enc_block_n910) );
  XNOR2X1 aes_core_enc_block_U826 ( .A(aes_core_round_key[36]), .B(Din[36]), 
        .Y(aes_core_enc_block_n909) );
  OAI221X1 aes_core_enc_block_U825 ( .A0(aes_core_enc_block_n909), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1350), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n910), .Y(
        aes_core_enc_block_n1301) );
  XNOR2X1 aes_core_enc_block_U824 ( .A(aes_core_round_key[12]), .B(
        aes_core_enc_block_n1368), .Y(aes_core_enc_block_n1095) );
  AOI222X1 aes_core_enc_block_U823 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[12]), .B0(aes_core_enc_block_n60), .B1(
        aes_core_enc_block_n1095), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1096), .Y(aes_core_enc_block_n1094) );
  XNOR2X1 aes_core_enc_block_U822 ( .A(aes_core_round_key[12]), .B(Din[12]), 
        .Y(aes_core_enc_block_n1093) );
  OAI221X1 aes_core_enc_block_U821 ( .A0(aes_core_enc_block_n1093), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1351), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1094), .Y(
        aes_core_enc_block_n1325) );
  XNOR2X1 aes_core_enc_block_U820 ( .A(aes_core_round_key[68]), .B(
        aes_core_enc_block_n1367), .Y(aes_core_enc_block_n670) );
  AOI222X1 aes_core_enc_block_U819 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[4]), .B0(aes_core_enc_block_n46), .B1(
        aes_core_enc_block_n670), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n671), .Y(aes_core_enc_block_n669) );
  XNOR2X1 aes_core_enc_block_U818 ( .A(aes_core_round_key[68]), .B(Din[68]), 
        .Y(aes_core_enc_block_n668) );
  OAI221X1 aes_core_enc_block_U817 ( .A0(aes_core_enc_block_n668), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1352), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n669), .Y(
        aes_core_enc_block_n1269) );
  XNOR2X1 aes_core_enc_block_U816 ( .A(aes_core_round_key[46]), .B(
        aes_core_enc_block_n196), .Y(aes_core_enc_block_n844) );
  AOI222X1 aes_core_enc_block_U815 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[14]), .B0(aes_core_enc_block_n52), .B1(
        aes_core_enc_block_n844), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n845), .Y(aes_core_enc_block_n843) );
  XNOR2X1 aes_core_enc_block_U814 ( .A(aes_core_round_key[46]), .B(Din[46]), 
        .Y(aes_core_enc_block_n842) );
  OAI221X1 aes_core_enc_block_U813 ( .A0(aes_core_enc_block_n842), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1356), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n843), .Y(
        aes_core_enc_block_n1291) );
  XNOR2X1 aes_core_enc_block_U812 ( .A(aes_core_round_key[70]), .B(
        aes_core_enc_block_n1357), .Y(aes_core_enc_block_n656) );
  AOI222X1 aes_core_enc_block_U811 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[6]), .B0(aes_core_enc_block_n45), .B1(
        aes_core_enc_block_n656), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n657), .Y(aes_core_enc_block_n655) );
  XNOR2X1 aes_core_enc_block_U810 ( .A(aes_core_round_key[70]), .B(Din[70]), 
        .Y(aes_core_enc_block_n654) );
  OAI221X1 aes_core_enc_block_U809 ( .A0(aes_core_enc_block_n654), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1358), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n655), .Y(
        aes_core_enc_block_n1267) );
  XNOR2X1 aes_core_enc_block_U808 ( .A(aes_core_round_key[84]), .B(
        aes_core_enc_block_n1401), .Y(aes_core_enc_block_n560) );
  AOI222X1 aes_core_enc_block_U807 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[20]), .B0(aes_core_enc_block_n40), .B1(
        aes_core_enc_block_n560), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n561), .Y(aes_core_enc_block_n559) );
  XNOR2X1 aes_core_enc_block_U806 ( .A(aes_core_round_key[84]), .B(Din[84]), 
        .Y(aes_core_enc_block_n558) );
  OAI221X1 aes_core_enc_block_U805 ( .A0(aes_core_enc_block_n558), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1366), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n559), .Y(
        aes_core_enc_block_n1253) );
  XNOR2X1 aes_core_enc_block_U804 ( .A(aes_core_round_key[76]), .B(
        aes_core_enc_block_n1351), .Y(aes_core_enc_block_n615) );
  AOI222X1 aes_core_enc_block_U803 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[12]), .B0(aes_core_enc_block_n42), .B1(
        aes_core_enc_block_n615), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n616), .Y(aes_core_enc_block_n614) );
  XNOR2X1 aes_core_enc_block_U802 ( .A(aes_core_round_key[76]), .B(Din[76]), 
        .Y(aes_core_enc_block_n613) );
  OAI221X1 aes_core_enc_block_U801 ( .A0(aes_core_enc_block_n613), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1368), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n614), .Y(
        aes_core_enc_block_n1261) );
  XNOR2X1 aes_core_enc_block_U800 ( .A(aes_core_round_key[78]), .B(
        aes_core_enc_block_n1381), .Y(aes_core_enc_block_n603) );
  AOI222X1 aes_core_enc_block_U799 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[14]), .B0(aes_core_enc_block_n42), .B1(
        aes_core_enc_block_n603), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n604), .Y(aes_core_enc_block_n602) );
  XNOR2X1 aes_core_enc_block_U798 ( .A(aes_core_round_key[78]), .B(Din[78]), 
        .Y(aes_core_enc_block_n601) );
  OAI221X1 aes_core_enc_block_U797 ( .A0(aes_core_enc_block_n601), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1370), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n602), .Y(
        aes_core_enc_block_n1259) );
  XNOR2X1 aes_core_enc_block_U796 ( .A(aes_core_round_key[44]), .B(
        aes_core_enc_block_n1349), .Y(aes_core_enc_block_n856) );
  AOI222X1 aes_core_enc_block_U795 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[12]), .B0(aes_core_enc_block_n53), .B1(
        aes_core_enc_block_n856), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n857), .Y(aes_core_enc_block_n855) );
  XNOR2X1 aes_core_enc_block_U794 ( .A(aes_core_round_key[44]), .B(Din[44]), 
        .Y(aes_core_enc_block_n854) );
  OAI221X1 aes_core_enc_block_U793 ( .A0(aes_core_enc_block_n854), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1377), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n855), .Y(
        aes_core_enc_block_n1293) );
  XNOR2X1 aes_core_enc_block_U792 ( .A(aes_core_round_key[14]), .B(
        aes_core_enc_block_n1370), .Y(aes_core_enc_block_n1083) );
  AOI222X1 aes_core_enc_block_U791 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[14]), .B0(aes_core_enc_block_n60), .B1(
        aes_core_enc_block_n1083), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1084), .Y(aes_core_enc_block_n1082) );
  XNOR2X1 aes_core_enc_block_U790 ( .A(aes_core_round_key[14]), .B(Din[14]), 
        .Y(aes_core_enc_block_n1081) );
  OAI221X1 aes_core_enc_block_U789 ( .A0(aes_core_enc_block_n1081), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1381), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1082), .Y(
        aes_core_enc_block_n1323) );
  XNOR2X1 aes_core_enc_block_U788 ( .A(aes_core_round_key[20]), .B(
        aes_core_enc_block_n1388), .Y(aes_core_enc_block_n1040) );
  AOI222X1 aes_core_enc_block_U787 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[20]), .B0(aes_core_enc_block_n58), .B1(
        aes_core_enc_block_n1040), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n1041), .Y(aes_core_enc_block_n1039) );
  XNOR2X1 aes_core_enc_block_U786 ( .A(aes_core_round_key[20]), .B(Din[20]), 
        .Y(aes_core_enc_block_n1038) );
  OAI221X1 aes_core_enc_block_U785 ( .A0(aes_core_enc_block_n1038), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1390), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1039), .Y(
        aes_core_enc_block_n1317) );
  XNOR2X1 aes_core_enc_block_U784 ( .A(aes_core_round_key[52]), .B(
        aes_core_enc_block_n1390), .Y(aes_core_enc_block_n801) );
  AOI222X1 aes_core_enc_block_U783 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[20]), .B0(aes_core_enc_block_n50), .B1(
        aes_core_enc_block_n801), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n802), .Y(aes_core_enc_block_n800) );
  XNOR2X1 aes_core_enc_block_U782 ( .A(aes_core_round_key[52]), .B(Din[52]), 
        .Y(aes_core_enc_block_n799) );
  OAI221X1 aes_core_enc_block_U781 ( .A0(aes_core_enc_block_n799), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1401), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n800), .Y(
        aes_core_enc_block_n1285) );
  XNOR2X1 aes_core_enc_block_U780 ( .A(aes_core_round_key[22]), .B(
        aes_core_enc_block_n1410), .Y(aes_core_enc_block_n1026) );
  AOI222X1 aes_core_enc_block_U779 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[22]), .B0(aes_core_enc_block_n57), .B1(
        aes_core_enc_block_n1026), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n1027), .Y(aes_core_enc_block_n1025) );
  XNOR2X1 aes_core_enc_block_U778 ( .A(aes_core_round_key[22]), .B(Din[22]), 
        .Y(aes_core_enc_block_n1024) );
  OAI221X1 aes_core_enc_block_U777 ( .A0(aes_core_enc_block_n1024), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1411), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1025), .Y(
        aes_core_enc_block_n1315) );
  XNOR2X1 aes_core_enc_block_U776 ( .A(aes_core_round_key[54]), .B(
        aes_core_enc_block_n1411), .Y(aes_core_enc_block_n787) );
  AOI222X1 aes_core_enc_block_U775 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[22]), .B0(aes_core_enc_block_n49), .B1(
        aes_core_enc_block_n787), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n788), .Y(aes_core_enc_block_n786) );
  XNOR2X1 aes_core_enc_block_U774 ( .A(aes_core_round_key[54]), .B(Din[54]), 
        .Y(aes_core_enc_block_n785) );
  OAI221X1 aes_core_enc_block_U773 ( .A0(aes_core_enc_block_n785), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1412), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n786), .Y(
        aes_core_enc_block_n1283) );
  XNOR2X1 aes_core_enc_block_U772 ( .A(aes_core_round_key[86]), .B(
        aes_core_enc_block_n1412), .Y(aes_core_enc_block_n546) );
  AOI222X1 aes_core_enc_block_U771 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[22]), .B0(aes_core_enc_block_n38), .B1(
        aes_core_enc_block_n546), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n547), .Y(aes_core_enc_block_n545) );
  XNOR2X1 aes_core_enc_block_U770 ( .A(aes_core_round_key[86]), .B(Din[86]), 
        .Y(aes_core_enc_block_n544) );
  OAI221X1 aes_core_enc_block_U769 ( .A0(aes_core_enc_block_n544), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1414), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n545), .Y(
        aes_core_enc_block_n1251) );
  XNOR2X1 aes_core_enc_block_U768 ( .A(aes_core_round_key[65]), .B(
        aes_core_enc_block_n1207), .Y(aes_core_enc_block_n693) );
  AOI222X1 aes_core_enc_block_U767 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[1]), .B0(aes_core_enc_block_n47), .B1(
        aes_core_enc_block_n693), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n694), .Y(aes_core_enc_block_n692) );
  XNOR2X1 aes_core_enc_block_U766 ( .A(aes_core_round_key[65]), .B(Din[65]), 
        .Y(aes_core_enc_block_n691) );
  OAI221X1 aes_core_enc_block_U765 ( .A0(aes_core_enc_block_n691), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n188), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n692), .Y(
        aes_core_enc_block_n1272) );
  XNOR2X1 aes_core_enc_block_U764 ( .A(aes_core_round_key[41]), .B(
        aes_core_enc_block_n1436), .Y(aes_core_enc_block_n877) );
  AOI222X1 aes_core_enc_block_U763 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[9]), .B0(aes_core_enc_block_n54), .B1(
        aes_core_enc_block_n877), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n878), .Y(aes_core_enc_block_n876) );
  XNOR2X1 aes_core_enc_block_U762 ( .A(aes_core_round_key[41]), .B(Din[41]), 
        .Y(aes_core_enc_block_n875) );
  OAI221X1 aes_core_enc_block_U761 ( .A0(aes_core_enc_block_n875), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1363), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n876), .Y(
        aes_core_enc_block_n1296) );
  XNOR2X1 aes_core_enc_block_U760 ( .A(aes_core_round_key[9]), .B(
        aes_core_enc_block_n1437), .Y(aes_core_enc_block_n1116) );
  AOI222X1 aes_core_enc_block_U759 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[9]), .B0(aes_core_enc_block_n62), .B1(
        aes_core_enc_block_n1116), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1117), .Y(aes_core_enc_block_n1115) );
  XNOR2X1 aes_core_enc_block_U758 ( .A(aes_core_round_key[9]), .B(Din[9]), .Y(
        aes_core_enc_block_n1114) );
  OAI221X1 aes_core_enc_block_U757 ( .A0(aes_core_enc_block_n1114), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1373), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1115), .Y(
        aes_core_enc_block_n1328) );
  XNOR2X1 aes_core_enc_block_U756 ( .A(aes_core_round_key[1]), .B(
        aes_core_enc_block_n1456), .Y(aes_core_enc_block_n1173) );
  AOI222X1 aes_core_enc_block_U755 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[1]), .B0(aes_core_enc_block_n64), .B1(
        aes_core_enc_block_n1173), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n1174), .Y(aes_core_enc_block_n1172) );
  XNOR2X1 aes_core_enc_block_U754 ( .A(aes_core_round_key[1]), .B(Din[1]), .Y(
        aes_core_enc_block_n1171) );
  OAI221X1 aes_core_enc_block_U753 ( .A0(aes_core_enc_block_n1171), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1397), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1172), .Y(
        aes_core_enc_block_n1336) );
  XNOR2X1 aes_core_enc_block_U752 ( .A(aes_core_round_key[73]), .B(
        aes_core_enc_block_n1373), .Y(aes_core_enc_block_n636) );
  AOI222X1 aes_core_enc_block_U751 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[9]), .B0(aes_core_enc_block_n43), .B1(
        aes_core_enc_block_n636), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n637), .Y(aes_core_enc_block_n635) );
  XNOR2X1 aes_core_enc_block_U750 ( .A(aes_core_round_key[73]), .B(Din[73]), 
        .Y(aes_core_enc_block_n634) );
  OAI221X1 aes_core_enc_block_U749 ( .A0(aes_core_enc_block_n634), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1437), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n635), .Y(
        aes_core_enc_block_n1264) );
  XNOR2X1 aes_core_enc_block_U748 ( .A(aes_core_round_key[33]), .B(
        aes_core_enc_block_n188), .Y(aes_core_enc_block_n934) );
  AOI222X1 aes_core_enc_block_U747 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[1]), .B0(aes_core_enc_block_n57), .B1(
        aes_core_enc_block_n934), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n935), .Y(aes_core_enc_block_n933) );
  XNOR2X1 aes_core_enc_block_U746 ( .A(aes_core_round_key[33]), .B(Din[33]), 
        .Y(aes_core_enc_block_n932) );
  OAI221X1 aes_core_enc_block_U745 ( .A0(aes_core_enc_block_n932), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1456), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n933), .Y(
        aes_core_enc_block_n1304) );
  XNOR2X1 aes_core_enc_block_U744 ( .A(aes_core_round_key[42]), .B(
        aes_core_enc_block_n1364), .Y(aes_core_enc_block_n871) );
  AOI222X1 aes_core_enc_block_U743 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[10]), .B0(aes_core_enc_block_n52), .B1(
        aes_core_enc_block_n871), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n872), .Y(aes_core_enc_block_n870) );
  XNOR2X1 aes_core_enc_block_U742 ( .A(aes_core_round_key[42]), .B(Din[42]), 
        .Y(aes_core_enc_block_n869) );
  OAI221X1 aes_core_enc_block_U741 ( .A0(aes_core_enc_block_n869), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n189), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n870), .Y(
        aes_core_enc_block_n1295) );
  XNOR2X1 aes_core_enc_block_U740 ( .A(aes_core_round_key[66]), .B(
        aes_core_enc_block_n1398), .Y(aes_core_enc_block_n686) );
  AOI222X1 aes_core_enc_block_U739 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[2]), .B0(aes_core_enc_block_n47), .B1(
        aes_core_enc_block_n686), .C0(aes_core_enc_block_n117), .C1(
        aes_core_enc_block_n687), .Y(aes_core_enc_block_n685) );
  XNOR2X1 aes_core_enc_block_U738 ( .A(aes_core_round_key[66]), .B(Din[66]), 
        .Y(aes_core_enc_block_n684) );
  OAI221X1 aes_core_enc_block_U737 ( .A0(aes_core_enc_block_n684), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1347), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n685), .Y(
        aes_core_enc_block_n1271) );
  XNOR2X1 aes_core_enc_block_U736 ( .A(aes_core_round_key[43]), .B(
        aes_core_enc_block_n190), .Y(aes_core_enc_block_n864) );
  AOI222X1 aes_core_enc_block_U735 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[11]), .B0(aes_core_enc_block_n52), .B1(
        aes_core_enc_block_n864), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n865), .Y(aes_core_enc_block_n863) );
  XNOR2X1 aes_core_enc_block_U734 ( .A(aes_core_round_key[43]), .B(Din[43]), 
        .Y(aes_core_enc_block_n862) );
  OAI221X1 aes_core_enc_block_U733 ( .A0(aes_core_enc_block_n862), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1348), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n863), .Y(
        aes_core_enc_block_n1294) );
  XNOR2X1 aes_core_enc_block_U732 ( .A(aes_core_round_key[74]), .B(
        aes_core_enc_block_n1458), .Y(aes_core_enc_block_n630) );
  AOI222X1 aes_core_enc_block_U731 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[10]), .B0(aes_core_enc_block_n43), .B1(
        aes_core_enc_block_n630), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n631), .Y(aes_core_enc_block_n629) );
  XNOR2X1 aes_core_enc_block_U730 ( .A(aes_core_round_key[74]), .B(Din[74]), 
        .Y(aes_core_enc_block_n628) );
  OAI221X1 aes_core_enc_block_U729 ( .A0(aes_core_enc_block_n628), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1374), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n629), .Y(
        aes_core_enc_block_n1263) );
  XNOR2X1 aes_core_enc_block_U728 ( .A(aes_core_round_key[11]), .B(
        aes_core_enc_block_n1399), .Y(aes_core_enc_block_n1103) );
  AOI222X1 aes_core_enc_block_U727 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[11]), .B0(aes_core_enc_block_n61), .B1(
        aes_core_enc_block_n1103), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1104), .Y(aes_core_enc_block_n1102) );
  XNOR2X1 aes_core_enc_block_U726 ( .A(aes_core_round_key[11]), .B(Din[11]), 
        .Y(aes_core_enc_block_n1101) );
  OAI221X1 aes_core_enc_block_U725 ( .A0(aes_core_enc_block_n1101), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1375), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1102), .Y(
        aes_core_enc_block_n1326) );
  XNOR2X1 aes_core_enc_block_U724 ( .A(aes_core_round_key[75]), .B(
        aes_core_enc_block_n1375), .Y(aes_core_enc_block_n623) );
  AOI222X1 aes_core_enc_block_U723 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[11]), .B0(aes_core_enc_block_n43), .B1(
        aes_core_enc_block_n623), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n624), .Y(aes_core_enc_block_n622) );
  XNOR2X1 aes_core_enc_block_U722 ( .A(aes_core_round_key[75]), .B(Din[75]), 
        .Y(aes_core_enc_block_n621) );
  OAI221X1 aes_core_enc_block_U721 ( .A0(aes_core_enc_block_n621), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1399), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n622), .Y(
        aes_core_enc_block_n1262) );
  XNOR2X1 aes_core_enc_block_U720 ( .A(aes_core_round_key[50]), .B(
        aes_core_enc_block_n1448), .Y(aes_core_enc_block_n817) );
  AOI222X1 aes_core_enc_block_U719 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[18]), .B0(aes_core_enc_block_n51), .B1(
        aes_core_enc_block_n817), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n818), .Y(aes_core_enc_block_n816) );
  XNOR2X1 aes_core_enc_block_U718 ( .A(aes_core_round_key[50]), .B(Din[50]), 
        .Y(aes_core_enc_block_n815) );
  OAI221X1 aes_core_enc_block_U717 ( .A0(aes_core_enc_block_n815), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1442), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n816), .Y(
        aes_core_enc_block_n1287) );
  XNOR2X1 aes_core_enc_block_U716 ( .A(aes_core_round_key[82]), .B(
        aes_core_enc_block_n1442), .Y(aes_core_enc_block_n576) );
  AOI222X1 aes_core_enc_block_U715 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[18]), .B0(aes_core_enc_block_n41), .B1(
        aes_core_enc_block_n576), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n577), .Y(aes_core_enc_block_n575) );
  XNOR2X1 aes_core_enc_block_U714 ( .A(aes_core_round_key[82]), .B(Din[82]), 
        .Y(aes_core_enc_block_n574) );
  OAI221X1 aes_core_enc_block_U713 ( .A0(aes_core_enc_block_n574), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1444), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n575), .Y(
        aes_core_enc_block_n1255) );
  XNOR2X1 aes_core_enc_block_U712 ( .A(aes_core_round_key[18]), .B(
        aes_core_enc_block_n1446), .Y(aes_core_enc_block_n1056) );
  AOI222X1 aes_core_enc_block_U711 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[18]), .B0(aes_core_enc_block_n59), .B1(
        aes_core_enc_block_n1056), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n1057), .Y(aes_core_enc_block_n1055) );
  XNOR2X1 aes_core_enc_block_U710 ( .A(aes_core_round_key[18]), .B(Din[18]), 
        .Y(aes_core_enc_block_n1054) );
  OAI221X1 aes_core_enc_block_U709 ( .A0(aes_core_enc_block_n1054), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1448), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1055), .Y(
        aes_core_enc_block_n1319) );
  XNOR2X1 aes_core_enc_block_U708 ( .A(aes_core_round_key[34]), .B(
        aes_core_enc_block_n1347), .Y(aes_core_enc_block_n927) );
  AOI222X1 aes_core_enc_block_U707 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[2]), .B0(aes_core_enc_block_n56), .B1(
        aes_core_enc_block_n927), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n928), .Y(aes_core_enc_block_n926) );
  XNOR2X1 aes_core_enc_block_U706 ( .A(aes_core_round_key[34]), .B(Din[34]), 
        .Y(aes_core_enc_block_n925) );
  OAI221X1 aes_core_enc_block_U705 ( .A0(aes_core_enc_block_n925), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1454), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n926), .Y(
        aes_core_enc_block_n1303) );
  XNOR2X1 aes_core_enc_block_U704 ( .A(aes_core_round_key[2]), .B(
        aes_core_enc_block_n1454), .Y(aes_core_enc_block_n1166) );
  AOI222X1 aes_core_enc_block_U703 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[2]), .B0(aes_core_enc_block_n64), .B1(
        aes_core_enc_block_n1166), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1167), .Y(aes_core_enc_block_n1165) );
  XNOR2X1 aes_core_enc_block_U702 ( .A(aes_core_round_key[2]), .B(Din[2]), .Y(
        aes_core_enc_block_n1164) );
  OAI221X1 aes_core_enc_block_U701 ( .A0(aes_core_enc_block_n1164), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1457), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1165), .Y(
        aes_core_enc_block_n1335) );
  XNOR2X1 aes_core_enc_block_U700 ( .A(aes_core_round_key[10]), .B(
        aes_core_enc_block_n1374), .Y(aes_core_enc_block_n1110) );
  AOI222X1 aes_core_enc_block_U699 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[10]), .B0(aes_core_enc_block_n61), .B1(
        aes_core_enc_block_n1110), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1111), .Y(aes_core_enc_block_n1109) );
  XNOR2X1 aes_core_enc_block_U698 ( .A(aes_core_round_key[10]), .B(Din[10]), 
        .Y(aes_core_enc_block_n1108) );
  OAI221X1 aes_core_enc_block_U697 ( .A0(aes_core_enc_block_n1108), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1458), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1109), .Y(
        aes_core_enc_block_n1327) );
  XNOR2X1 aes_core_enc_block_U696 ( .A(aes_core_round_key[109]), .B(
        aes_core_enc_block_n1353), .Y(aes_core_enc_block_n377) );
  AOI222X1 aes_core_enc_block_U695 ( .A0(aes_core_new_sboxw[13]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n33), .B1(
        aes_core_enc_block_n377), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n378), .Y(aes_core_enc_block_n376) );
  XNOR2X1 aes_core_enc_block_U694 ( .A(aes_core_round_key[109]), .B(Din[109]), 
        .Y(aes_core_enc_block_n375) );
  OAI221X1 aes_core_enc_block_U693 ( .A0(aes_core_enc_block_n375), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n193), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n376), .Y(
        aes_core_enc_block_n1229) );
  XNOR2X1 aes_core_enc_block_U692 ( .A(aes_core_round_key[111]), .B(
        aes_core_enc_block_n1359), .Y(aes_core_enc_block_n365) );
  AOI222X1 aes_core_enc_block_U691 ( .A0(aes_core_new_sboxw[15]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n32), .B1(
        aes_core_enc_block_n365), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n366), .Y(aes_core_enc_block_n364) );
  XNOR2X1 aes_core_enc_block_U690 ( .A(aes_core_round_key[111]), .B(Din[111]), 
        .Y(aes_core_enc_block_n363) );
  OAI221X1 aes_core_enc_block_U689 ( .A0(aes_core_enc_block_n363), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n467), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n364), .Y(
        aes_core_enc_block_n1227) );
  XNOR2X1 aes_core_enc_block_U688 ( .A(aes_core_round_key[37]), .B(
        aes_core_enc_block_n1355), .Y(aes_core_enc_block_n904) );
  AOI222X1 aes_core_enc_block_U687 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[5]), .B0(aes_core_enc_block_n55), .B1(
        aes_core_enc_block_n904), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n905), .Y(aes_core_enc_block_n903) );
  XNOR2X1 aes_core_enc_block_U686 ( .A(aes_core_round_key[37]), .B(Din[37]), 
        .Y(aes_core_enc_block_n902) );
  OAI221X1 aes_core_enc_block_U685 ( .A0(aes_core_enc_block_n902), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n194), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n903), .Y(
        aes_core_enc_block_n1300) );
  XNOR2X1 aes_core_enc_block_U684 ( .A(aes_core_round_key[5]), .B(
        aes_core_enc_block_n194), .Y(aes_core_enc_block_n1143) );
  AOI222X1 aes_core_enc_block_U683 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[5]), .B0(aes_core_enc_block_n63), .B1(
        aes_core_enc_block_n1143), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1144), .Y(aes_core_enc_block_n1142) );
  XNOR2X1 aes_core_enc_block_U682 ( .A(aes_core_round_key[5]), .B(Din[5]), .Y(
        aes_core_enc_block_n1141) );
  OAI221X1 aes_core_enc_block_U681 ( .A0(aes_core_enc_block_n1141), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n195), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1142), .Y(
        aes_core_enc_block_n1332) );
  XNOR2X1 aes_core_enc_block_U680 ( .A(aes_core_round_key[45]), .B(
        aes_core_enc_block_n193), .Y(aes_core_enc_block_n850) );
  AOI222X1 aes_core_enc_block_U679 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[13]), .B0(aes_core_enc_block_n53), .B1(
        aes_core_enc_block_n850), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n851), .Y(aes_core_enc_block_n849) );
  XNOR2X1 aes_core_enc_block_U678 ( .A(aes_core_round_key[45]), .B(Din[45]), 
        .Y(aes_core_enc_block_n848) );
  OAI221X1 aes_core_enc_block_U677 ( .A0(aes_core_enc_block_n848), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1353), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n849), .Y(
        aes_core_enc_block_n1292) );
  XNOR2X1 aes_core_enc_block_U676 ( .A(aes_core_round_key[69]), .B(
        aes_core_enc_block_n1354), .Y(aes_core_enc_block_n663) );
  AOI222X1 aes_core_enc_block_U675 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[5]), .B0(aes_core_enc_block_n45), .B1(
        aes_core_enc_block_n663), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n664), .Y(aes_core_enc_block_n662) );
  XNOR2X1 aes_core_enc_block_U674 ( .A(aes_core_round_key[69]), .B(Din[69]), 
        .Y(aes_core_enc_block_n661) );
  OAI221X1 aes_core_enc_block_U673 ( .A0(aes_core_enc_block_n661), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1355), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n662), .Y(
        aes_core_enc_block_n1268) );
  XNOR2X1 aes_core_enc_block_U672 ( .A(aes_core_round_key[47]), .B(
        aes_core_enc_block_n467), .Y(aes_core_enc_block_n838) );
  AOI222X1 aes_core_enc_block_U671 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[15]), .B0(aes_core_enc_block_n52), .B1(
        aes_core_enc_block_n838), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n839), .Y(aes_core_enc_block_n837) );
  XNOR2X1 aes_core_enc_block_U670 ( .A(aes_core_round_key[47]), .B(Din[47]), 
        .Y(aes_core_enc_block_n836) );
  OAI221X1 aes_core_enc_block_U669 ( .A0(aes_core_enc_block_n836), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1359), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n837), .Y(
        aes_core_enc_block_n1290) );
  XNOR2X1 aes_core_enc_block_U668 ( .A(aes_core_round_key[13]), .B(
        aes_core_enc_block_n1404), .Y(aes_core_enc_block_n1089) );
  AOI222X1 aes_core_enc_block_U667 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[13]), .B0(aes_core_enc_block_n61), .B1(
        aes_core_enc_block_n1089), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1090), .Y(aes_core_enc_block_n1088) );
  XNOR2X1 aes_core_enc_block_U666 ( .A(aes_core_round_key[13]), .B(Din[13]), 
        .Y(aes_core_enc_block_n1087) );
  OAI221X1 aes_core_enc_block_U665 ( .A0(aes_core_enc_block_n1087), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1369), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1088), .Y(
        aes_core_enc_block_n1324) );
  XNOR2X1 aes_core_enc_block_U664 ( .A(aes_core_round_key[15]), .B(
        aes_core_enc_block_n1382), .Y(aes_core_enc_block_n1077) );
  AOI222X1 aes_core_enc_block_U663 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[15]), .B0(aes_core_enc_block_n60), .B1(
        aes_core_enc_block_n1077), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1078), .Y(aes_core_enc_block_n1076) );
  XNOR2X1 aes_core_enc_block_U662 ( .A(aes_core_round_key[15]), .B(Din[15]), 
        .Y(aes_core_enc_block_n1075) );
  OAI221X1 aes_core_enc_block_U661 ( .A0(aes_core_enc_block_n1075), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1371), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1076), .Y(
        aes_core_enc_block_n1322) );
  XNOR2X1 aes_core_enc_block_U660 ( .A(aes_core_round_key[79]), .B(
        aes_core_enc_block_n1371), .Y(aes_core_enc_block_n597) );
  AOI222X1 aes_core_enc_block_U659 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[15]), .B0(aes_core_enc_block_n41), .B1(
        aes_core_enc_block_n597), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n598), .Y(aes_core_enc_block_n596) );
  XNOR2X1 aes_core_enc_block_U658 ( .A(aes_core_round_key[79]), .B(Din[79]), 
        .Y(aes_core_enc_block_n595) );
  OAI221X1 aes_core_enc_block_U657 ( .A0(aes_core_enc_block_n595), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1382), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n596), .Y(
        aes_core_enc_block_n1258) );
  XNOR2X1 aes_core_enc_block_U656 ( .A(aes_core_round_key[77]), .B(
        aes_core_enc_block_n1369), .Y(aes_core_enc_block_n609) );
  AOI222X1 aes_core_enc_block_U655 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[13]), .B0(aes_core_enc_block_n42), .B1(
        aes_core_enc_block_n609), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n610), .Y(aes_core_enc_block_n608) );
  XNOR2X1 aes_core_enc_block_U654 ( .A(aes_core_round_key[77]), .B(Din[77]), 
        .Y(aes_core_enc_block_n607) );
  OAI221X1 aes_core_enc_block_U653 ( .A0(aes_core_enc_block_n607), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1404), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n608), .Y(
        aes_core_enc_block_n1260) );
  AOI22X1 aes_core_enc_block_U652 ( .A0(Dout[29]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[61]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n208) );
  OAI221X1 aes_core_enc_block_U651 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1403), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1408), .C0(aes_core_enc_block_n208), .Y(
        aes_core_enc_sboxw[29]) );
  AOI22X1 aes_core_enc_block_U650 ( .A0(Dout[26]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[58]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n211) );
  OAI221X1 aes_core_enc_block_U649 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1443), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1445), .C0(aes_core_enc_block_n211), .Y(
        aes_core_enc_sboxw[26]) );
  XNOR2X1 aes_core_enc_block_U648 ( .A(aes_core_round_key[115]), .B(
        aes_core_enc_block_n1386), .Y(aes_core_enc_block_n336) );
  AOI222X1 aes_core_enc_block_U647 ( .A0(aes_core_new_sboxw[19]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n30), .B1(
        aes_core_enc_block_n336), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n337), .Y(aes_core_enc_block_n335) );
  XNOR2X1 aes_core_enc_block_U646 ( .A(aes_core_round_key[115]), .B(Din[115]), 
        .Y(aes_core_enc_block_n334) );
  OAI221X1 aes_core_enc_block_U645 ( .A0(aes_core_enc_block_n334), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1450), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n335), .Y(
        aes_core_enc_block_n1223) );
  OAI2BB2X1 aes_core_enc_block_U644 ( .B0(aes_core_enc_block_n1394), .B1(
        aes_core_enc_block_n26), .A0N(aes_core_enc_block_n112), .A1N(Din[63]), 
        .Y(aes_core_enc_block_n712) );
  XOR2X1 aes_core_enc_block_U643 ( .A(aes_core_enc_block_n714), .B(
        aes_core_enc_block_n715), .Y(aes_core_enc_block_n711) );
  AOI222X1 aes_core_enc_block_U642 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n711), .B0(aes_core_enc_block_n712), .B1(
        aes_core_enc_block_n148), .C0(aes_core_round_key[63]), .C1(
        aes_core_enc_block_n713), .Y(aes_core_enc_block_n710) );
  OAI221X1 aes_core_enc_block_U641 ( .A0(aes_core_enc_block_n159), .A1(
        aes_core_enc_block_n2), .B0(aes_core_enc_block_n1394), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n710), .Y(
        aes_core_enc_block_n1274) );
  OAI2BB2X1 aes_core_enc_block_U640 ( .B0(aes_core_enc_block_n1383), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n114), .A1N(Din[31]), 
        .Y(aes_core_enc_block_n951) );
  XOR2X1 aes_core_enc_block_U639 ( .A(aes_core_enc_block_n953), .B(
        aes_core_enc_block_n954), .Y(aes_core_enc_block_n950) );
  AOI222X1 aes_core_enc_block_U638 ( .A0(aes_core_enc_block_n121), .A1(
        aes_core_enc_block_n950), .B0(aes_core_enc_block_n951), .B1(
        aes_core_enc_block_n156), .C0(aes_core_round_key[31]), .C1(
        aes_core_enc_block_n952), .Y(aes_core_enc_block_n949) );
  OAI221X1 aes_core_enc_block_U637 ( .A0(aes_core_enc_block_n159), .A1(
        aes_core_enc_block_n4), .B0(aes_core_enc_block_n1383), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n949), .Y(
        aes_core_enc_block_n1306) );
  XNOR2X1 aes_core_enc_block_U636 ( .A(aes_core_round_key[87]), .B(
        aes_core_enc_block_n1416), .Y(aes_core_enc_block_n538) );
  AOI222X1 aes_core_enc_block_U635 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[23]), .B0(aes_core_enc_block_n39), .B1(
        aes_core_enc_block_n538), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n539), .Y(aes_core_enc_block_n537) );
  XNOR2X1 aes_core_enc_block_U634 ( .A(aes_core_round_key[87]), .B(Din[87]), 
        .Y(aes_core_enc_block_n536) );
  OAI221X1 aes_core_enc_block_U633 ( .A0(aes_core_enc_block_n536), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n1417), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n537), .Y(
        aes_core_enc_block_n1250) );
  XNOR2X1 aes_core_enc_block_U632 ( .A(aes_core_round_key[55]), .B(
        aes_core_enc_block_n1419), .Y(aes_core_enc_block_n779) );
  AOI222X1 aes_core_enc_block_U631 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[23]), .B0(aes_core_enc_block_n48), .B1(
        aes_core_enc_block_n779), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n780), .Y(aes_core_enc_block_n778) );
  XNOR2X1 aes_core_enc_block_U630 ( .A(aes_core_round_key[55]), .B(Din[55]), 
        .Y(aes_core_enc_block_n777) );
  OAI221X1 aes_core_enc_block_U629 ( .A0(aes_core_enc_block_n777), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1416), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n778), .Y(
        aes_core_enc_block_n1282) );
  XNOR2X1 aes_core_enc_block_U628 ( .A(aes_core_round_key[23]), .B(
        aes_core_enc_block_n1418), .Y(aes_core_enc_block_n1018) );
  AOI222X1 aes_core_enc_block_U627 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[23]), .B0(aes_core_enc_block_n57), .B1(
        aes_core_enc_block_n1018), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n1019), .Y(aes_core_enc_block_n1017) );
  XNOR2X1 aes_core_enc_block_U626 ( .A(aes_core_round_key[23]), .B(Din[23]), 
        .Y(aes_core_enc_block_n1016) );
  OAI221X1 aes_core_enc_block_U625 ( .A0(aes_core_enc_block_n1016), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1419), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1017), .Y(
        aes_core_enc_block_n1314) );
  OAI2BB2X1 aes_core_enc_block_U624 ( .B0(aes_core_enc_block_n1361), .B1(
        aes_core_enc_block_n25), .A0N(aes_core_enc_block_n108), .A1N(Din[95]), 
        .Y(aes_core_enc_block_n471) );
  XOR2X1 aes_core_enc_block_U623 ( .A(aes_core_enc_block_n473), .B(
        aes_core_enc_block_n474), .Y(aes_core_enc_block_n470) );
  AOI222X1 aes_core_enc_block_U622 ( .A0(aes_core_enc_block_n117), .A1(
        aes_core_enc_block_n470), .B0(aes_core_enc_block_n471), .B1(
        aes_core_enc_block_n140), .C0(aes_core_round_key[95]), .C1(
        aes_core_enc_block_n472), .Y(aes_core_enc_block_n469) );
  OAI221X1 aes_core_enc_block_U621 ( .A0(aes_core_enc_block_n159), .A1(
        aes_core_enc_block_n5), .B0(aes_core_enc_block_n1361), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n469), .Y(
        aes_core_enc_block_n1242) );
  OAI2BB2X1 aes_core_enc_block_U620 ( .B0(aes_core_enc_block_n1420), .B1(
        aes_core_enc_block_n24), .A0N(aes_core_enc_block_n112), .A1N(Din[127]), 
        .Y(aes_core_enc_block_n237) );
  XOR2X1 aes_core_enc_block_U619 ( .A(aes_core_enc_block_n241), .B(
        aes_core_enc_block_n242), .Y(aes_core_enc_block_n236) );
  AOI222X1 aes_core_enc_block_U618 ( .A0(aes_core_enc_block_n120), .A1(
        aes_core_enc_block_n236), .B0(aes_core_enc_block_n237), .B1(
        aes_core_enc_block_n132), .C0(aes_core_round_key[127]), .C1(
        aes_core_enc_block_n238), .Y(aes_core_enc_block_n234) );
  OAI221X1 aes_core_enc_block_U617 ( .A0(aes_core_enc_block_n3), .A1(
        aes_core_enc_block_n159), .B0(aes_core_enc_block_n1420), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n234), .Y(
        aes_core_enc_block_n1211) );
  XNOR2X1 aes_core_enc_block_U616 ( .A(aes_core_round_key[119]), .B(
        aes_core_enc_block_n1417), .Y(aes_core_enc_block_n306) );
  AOI222X1 aes_core_enc_block_U615 ( .A0(aes_core_new_sboxw[23]), .A1(
        aes_core_enc_block_n7), .B0(aes_core_enc_block_n50), .B1(
        aes_core_enc_block_n306), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n307), .Y(aes_core_enc_block_n305) );
  XNOR2X1 aes_core_enc_block_U614 ( .A(aes_core_round_key[119]), .B(Din[119]), 
        .Y(aes_core_enc_block_n304) );
  OAI221X1 aes_core_enc_block_U613 ( .A0(aes_core_enc_block_n304), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1418), .B1(
        aes_core_enc_block_n233), .C0(aes_core_enc_block_n305), .Y(
        aes_core_enc_block_n1219) );
  XNOR2X1 aes_core_enc_block_U612 ( .A(aes_core_round_key[35]), .B(
        aes_core_enc_block_n1376), .Y(aes_core_enc_block_n919) );
  AOI222X1 aes_core_enc_block_U611 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[3]), .B0(aes_core_enc_block_n56), .B1(
        aes_core_enc_block_n919), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n920), .Y(aes_core_enc_block_n918) );
  XNOR2X1 aes_core_enc_block_U610 ( .A(aes_core_round_key[35]), .B(Din[35]), 
        .Y(aes_core_enc_block_n917) );
  OAI221X1 aes_core_enc_block_U609 ( .A0(aes_core_enc_block_n917), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n191), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n918), .Y(
        aes_core_enc_block_n1302) );
  XNOR2X1 aes_core_enc_block_U608 ( .A(aes_core_round_key[51]), .B(
        aes_core_enc_block_n1400), .Y(aes_core_enc_block_n809) );
  AOI222X1 aes_core_enc_block_U607 ( .A0(aes_core_enc_block_n16), .A1(
        aes_core_new_sboxw[19]), .B0(aes_core_enc_block_n51), .B1(
        aes_core_enc_block_n809), .C0(aes_core_enc_block_n121), .C1(
        aes_core_enc_block_n810), .Y(aes_core_enc_block_n808) );
  XNOR2X1 aes_core_enc_block_U606 ( .A(aes_core_round_key[51]), .B(Din[51]), 
        .Y(aes_core_enc_block_n807) );
  OAI221X1 aes_core_enc_block_U605 ( .A0(aes_core_enc_block_n807), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1365), .B1(
        aes_core_enc_block_n709), .C0(aes_core_enc_block_n808), .Y(
        aes_core_enc_block_n1286) );
  XNOR2X1 aes_core_enc_block_U604 ( .A(aes_core_round_key[67]), .B(
        aes_core_enc_block_n1385), .Y(aes_core_enc_block_n678) );
  AOI222X1 aes_core_enc_block_U603 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[3]), .B0(aes_core_enc_block_n46), .B1(
        aes_core_enc_block_n678), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n679), .Y(aes_core_enc_block_n677) );
  XNOR2X1 aes_core_enc_block_U602 ( .A(aes_core_round_key[67]), .B(Din[67]), 
        .Y(aes_core_enc_block_n676) );
  OAI221X1 aes_core_enc_block_U601 ( .A0(aes_core_enc_block_n676), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1376), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n677), .Y(
        aes_core_enc_block_n1270) );
  XNOR2X1 aes_core_enc_block_U600 ( .A(aes_core_round_key[83]), .B(
        aes_core_enc_block_n1365), .Y(aes_core_enc_block_n568) );
  AOI222X1 aes_core_enc_block_U599 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[19]), .B0(aes_core_enc_block_n40), .B1(
        aes_core_enc_block_n568), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n569), .Y(aes_core_enc_block_n567) );
  XNOR2X1 aes_core_enc_block_U598 ( .A(aes_core_round_key[83]), .B(Din[83]), 
        .Y(aes_core_enc_block_n566) );
  OAI221X1 aes_core_enc_block_U597 ( .A0(aes_core_enc_block_n566), .A1(
        aes_core_enc_block_n101), .B0(aes_core_enc_block_n1386), .B1(
        aes_core_enc_block_n468), .C0(aes_core_enc_block_n567), .Y(
        aes_core_enc_block_n1254) );
  XNOR2X1 aes_core_enc_block_U596 ( .A(aes_core_round_key[19]), .B(
        aes_core_enc_block_n1450), .Y(aes_core_enc_block_n1048) );
  AOI222X1 aes_core_enc_block_U595 ( .A0(aes_core_enc_block_n12), .A1(
        aes_core_new_sboxw[19]), .B0(aes_core_enc_block_n59), .B1(
        aes_core_enc_block_n1048), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n1049), .Y(aes_core_enc_block_n1047) );
  XNOR2X1 aes_core_enc_block_U594 ( .A(aes_core_round_key[19]), .B(Din[19]), 
        .Y(aes_core_enc_block_n1046) );
  OAI221X1 aes_core_enc_block_U593 ( .A0(aes_core_enc_block_n1046), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1400), .B1(
        aes_core_enc_block_n948), .C0(aes_core_enc_block_n1047), .Y(
        aes_core_enc_block_n1318) );
  XNOR2X1 aes_core_enc_block_U592 ( .A(aes_core_round_key[3]), .B(
        aes_core_enc_block_n191), .Y(aes_core_enc_block_n1158) );
  AOI222X1 aes_core_enc_block_U591 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[3]), .B0(aes_core_enc_block_n64), .B1(
        aes_core_enc_block_n1158), .C0(aes_core_enc_block_n120), .C1(
        aes_core_enc_block_n1159), .Y(aes_core_enc_block_n1157) );
  XNOR2X1 aes_core_enc_block_U590 ( .A(aes_core_round_key[3]), .B(Din[3]), .Y(
        aes_core_enc_block_n1156) );
  OAI221X1 aes_core_enc_block_U589 ( .A0(aes_core_enc_block_n1156), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1455), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1157), .Y(
        aes_core_enc_block_n1334) );
  XNOR2X1 aes_core_enc_block_U588 ( .A(aes_core_round_key[103]), .B(
        aes_core_enc_block_n1384), .Y(aes_core_enc_block_n417) );
  AOI222X1 aes_core_enc_block_U587 ( .A0(aes_core_new_sboxw[7]), .A1(
        aes_core_enc_block_n8), .B0(aes_core_enc_block_n36), .B1(
        aes_core_enc_block_n417), .C0(aes_core_enc_block_n118), .C1(
        aes_core_enc_block_n418), .Y(aes_core_enc_block_n416) );
  XNOR2X1 aes_core_enc_block_U586 ( .A(aes_core_round_key[103]), .B(Din[103]), 
        .Y(aes_core_enc_block_n415) );
  OAI221X1 aes_core_enc_block_U585 ( .A0(aes_core_enc_block_n415), .A1(
        aes_core_enc_block_n104), .B0(aes_core_enc_block_n1360), .B1(
        aes_core_enc_block_n123), .C0(aes_core_enc_block_n416), .Y(
        aes_core_enc_block_n1235) );
  XNOR2X1 aes_core_enc_block_U584 ( .A(aes_core_round_key[39]), .B(
        aes_core_enc_block_n1415), .Y(aes_core_enc_block_n890) );
  AOI222X1 aes_core_enc_block_U583 ( .A0(aes_core_enc_block_n17), .A1(
        aes_core_new_sboxw[7]), .B0(aes_core_enc_block_n54), .B1(
        aes_core_enc_block_n890), .C0(aes_core_enc_block_n235), .C1(
        aes_core_enc_block_n891), .Y(aes_core_enc_block_n889) );
  XNOR2X1 aes_core_enc_block_U582 ( .A(aes_core_round_key[39]), .B(Din[39]), 
        .Y(aes_core_enc_block_n888) );
  OAI221X1 aes_core_enc_block_U581 ( .A0(aes_core_enc_block_n888), .A1(
        aes_core_enc_block_n103), .B0(aes_core_enc_block_n708), .B1(
        aes_core_enc_block_n20), .C0(aes_core_enc_block_n889), .Y(
        aes_core_enc_block_n1298) );
  XNOR2X1 aes_core_enc_block_U580 ( .A(aes_core_round_key[7]), .B(
        aes_core_enc_block_n708), .Y(aes_core_enc_block_n1129) );
  AOI222X1 aes_core_enc_block_U579 ( .A0(aes_core_enc_block_n13), .A1(
        aes_core_new_sboxw[7]), .B0(aes_core_enc_block_n62), .B1(
        aes_core_enc_block_n1129), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n1130), .Y(aes_core_enc_block_n1128) );
  XNOR2X1 aes_core_enc_block_U578 ( .A(aes_core_round_key[7]), .B(Din[7]), .Y(
        aes_core_enc_block_n1127) );
  OAI221X1 aes_core_enc_block_U577 ( .A0(aes_core_enc_block_n1127), .A1(
        aes_core_enc_block_n105), .B0(aes_core_enc_block_n1384), .B1(
        aes_core_enc_block_n18), .C0(aes_core_enc_block_n1128), .Y(
        aes_core_enc_block_n1330) );
  XNOR2X1 aes_core_enc_block_U576 ( .A(aes_core_round_key[71]), .B(
        aes_core_enc_block_n1360), .Y(aes_core_enc_block_n649) );
  AOI222X1 aes_core_enc_block_U575 ( .A0(aes_core_enc_block_n9), .A1(
        aes_core_new_sboxw[7]), .B0(aes_core_enc_block_n44), .B1(
        aes_core_enc_block_n649), .C0(aes_core_enc_block_n119), .C1(
        aes_core_enc_block_n650), .Y(aes_core_enc_block_n648) );
  XNOR2X1 aes_core_enc_block_U574 ( .A(aes_core_round_key[71]), .B(Din[71]), 
        .Y(aes_core_enc_block_n647) );
  OAI221X1 aes_core_enc_block_U573 ( .A0(aes_core_enc_block_n647), .A1(
        aes_core_enc_block_n102), .B0(aes_core_enc_block_n1415), .B1(
        aes_core_enc_block_n22), .C0(aes_core_enc_block_n648), .Y(
        aes_core_enc_block_n1266) );
  AOI22X1 aes_core_enc_block_U572 ( .A0(Dout[5]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[37]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n202) );
  OAI221X1 aes_core_enc_block_U571 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1355), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1354), .C0(aes_core_enc_block_n202), .Y(
        aes_core_enc_sboxw[5]) );
  AOI22X1 aes_core_enc_block_U570 ( .A0(Dout[21]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[53]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n216) );
  OAI221X1 aes_core_enc_block_U569 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1407), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1378), .C0(aes_core_enc_block_n216), .Y(
        aes_core_enc_sboxw[21]) );
  AOI22X1 aes_core_enc_block_U568 ( .A0(Dout[0]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[32]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n229) );
  OAI221X1 aes_core_enc_block_U567 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1362), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n187), .C0(aes_core_enc_block_n229), .Y(
        aes_core_enc_sboxw[0]) );
  AOI22X1 aes_core_enc_block_U566 ( .A0(Dout[1]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[33]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n218) );
  OAI221X1 aes_core_enc_block_U565 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n188), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1207), .C0(aes_core_enc_block_n218), .Y(
        aes_core_enc_sboxw[1]) );
  AOI22X1 aes_core_enc_block_U564 ( .A0(Dout[16]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[48]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n222) );
  OAI221X1 aes_core_enc_block_U563 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1430), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1424), .C0(aes_core_enc_block_n222), .Y(
        aes_core_enc_sboxw[16]) );
  AOI22X1 aes_core_enc_block_U562 ( .A0(Dout[17]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[49]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n221) );
  OAI221X1 aes_core_enc_block_U561 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1433), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1435), .C0(aes_core_enc_block_n221), .Y(
        aes_core_enc_sboxw[17]) );
  AOI22X1 aes_core_enc_block_U560 ( .A0(Dout[24]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[56]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n213) );
  OAI221X1 aes_core_enc_block_U559 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1429), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1421), .C0(aes_core_enc_block_n213), .Y(
        aes_core_enc_sboxw[24]) );
  AOI22X1 aes_core_enc_block_U558 ( .A0(Dout[25]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[57]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n212) );
  OAI221X1 aes_core_enc_block_U557 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1432), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1434), .C0(aes_core_enc_block_n212), .Y(
        aes_core_enc_sboxw[25]) );
  AOI22X1 aes_core_enc_block_U556 ( .A0(Dout[2]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[34]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n207) );
  AOI22X1 aes_core_enc_block_U555 ( .A0(Dout[9]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[41]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n198) );
  AOI22X1 aes_core_enc_block_U554 ( .A0(Dout[12]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[44]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n226) );
  AOI22X1 aes_core_enc_block_U553 ( .A0(Dout[8]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[40]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n199) );
  AOI22X1 aes_core_enc_block_U552 ( .A0(Dout[10]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[42]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n228) );
  AOI22X1 aes_core_enc_block_U551 ( .A0(Dout[18]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[50]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n220) );
  AOI22X1 aes_core_enc_block_U550 ( .A0(Dout[28]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[60]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n209) );
  AOI22X1 aes_core_enc_block_U549 ( .A0(Dout[13]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[45]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n225) );
  OAI221X1 aes_core_enc_block_U548 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1404), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n193), .C0(aes_core_enc_block_n225), .Y(
        aes_core_enc_sboxw[13]) );
  NOR2X1 aes_core_enc_block_U547 ( .A(aes_core_enc_block_enc_ctrl_reg[0]), .B(
        aes_core_enc_block_n180), .Y(aes_core_enc_block_n1195) );
  AOI22X1 aes_core_enc_block_U546 ( .A0(Dout[11]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[43]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n227) );
  OAI221X1 aes_core_enc_block_U545 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1399), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n190), .C0(aes_core_enc_block_n227), .Y(
        aes_core_enc_sboxw[11]) );
  AOI22X1 aes_core_enc_block_U544 ( .A0(Dout[27]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[59]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n210) );
  OAI221X1 aes_core_enc_block_U543 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1452), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1449), .C0(aes_core_enc_block_n210), .Y(
        aes_core_enc_sboxw[27]) );
  AOI22X1 aes_core_enc_block_U542 ( .A0(Dout[4]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[36]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n203) );
  AOI22X1 aes_core_enc_block_U541 ( .A0(Dout[20]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[52]), .B1(aes_core_enc_block_n15), .Y(aes_core_enc_block_n217) );
  AOI22X1 aes_core_enc_block_U540 ( .A0(Dout[3]), .A1(aes_core_enc_block_n11), 
        .B0(Dout[35]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n204) );
  AOI22X1 aes_core_enc_block_U539 ( .A0(Dout[19]), .A1(aes_core_enc_block_n10), 
        .B0(Dout[51]), .B1(aes_core_enc_block_n14), .Y(aes_core_enc_block_n219) );
  OAI221X1 aes_core_enc_block_U538 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1386), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1450), .C0(aes_core_enc_block_n219), .Y(
        aes_core_enc_sboxw[19]) );
  NOR2X1 aes_core_enc_block_U537 ( .A(aes_core_enc_block_n182), .B(
        aes_core_enc_block_n1203), .Y(aes_core_enc_block_n1200) );
  XOR2X1 aes_core_enc_block_U536 ( .A(aes_core_enc_block_n475), .B(
        aes_core_enc_block_n476), .Y(aes_core_enc_block_n474) );
  XOR2X1 aes_core_enc_block_U535 ( .A(aes_core_enc_block_n963), .B(
        aes_core_enc_block_n964), .Y(aes_core_enc_block_n962) );
  XOR2X1 aes_core_enc_block_U534 ( .A(aes_core_enc_block_n955), .B(
        aes_core_enc_block_n956), .Y(aes_core_enc_block_n954) );
  XOR2X1 aes_core_enc_block_U533 ( .A(aes_core_enc_block_n267), .B(
        aes_core_enc_block_n268), .Y(aes_core_enc_block_n266) );
  XOR2X1 aes_core_enc_block_U532 ( .A(aes_core_enc_block_n740), .B(
        aes_core_enc_block_n741), .Y(aes_core_enc_block_n739) );
  XOR2X1 aes_core_enc_block_U531 ( .A(aes_core_enc_block_n724), .B(
        aes_core_enc_block_n725), .Y(aes_core_enc_block_n723) );
  XOR2X1 aes_core_enc_block_U530 ( .A(aes_core_enc_block_n716), .B(
        aes_core_enc_block_n717), .Y(aes_core_enc_block_n715) );
  XOR2X1 aes_core_enc_block_U529 ( .A(aes_core_enc_block_n499), .B(
        aes_core_enc_block_n500), .Y(aes_core_enc_block_n498) );
  XOR2X1 aes_core_enc_block_U528 ( .A(aes_core_enc_block_n251), .B(
        aes_core_enc_block_n252), .Y(aes_core_enc_block_n250) );
  XOR2X1 aes_core_enc_block_U527 ( .A(aes_core_enc_block_n243), .B(
        aes_core_enc_block_n244), .Y(aes_core_enc_block_n242) );
  XOR2X1 aes_core_enc_block_U526 ( .A(aes_core_enc_block_n759), .B(
        aes_core_enc_block_n760), .Y(aes_core_enc_block_n758) );
  XOR2X1 aes_core_enc_block_U525 ( .A(aes_core_enc_block_n518), .B(
        aes_core_enc_block_n519), .Y(aes_core_enc_block_n517) );
  XOR2X1 aes_core_enc_block_U524 ( .A(aes_core_enc_block_n998), .B(
        aes_core_enc_block_n999), .Y(aes_core_enc_block_n997) );
  XOR2X1 aes_core_enc_block_U523 ( .A(aes_core_enc_block_n483), .B(
        aes_core_enc_block_n484), .Y(aes_core_enc_block_n482) );
  XOR2X1 aes_core_enc_block_U522 ( .A(aes_core_enc_block_n286), .B(
        aes_core_enc_block_n287), .Y(aes_core_enc_block_n285) );
  XOR2X1 aes_core_enc_block_U521 ( .A(aes_core_enc_block_n277), .B(
        aes_core_enc_block_n278), .Y(aes_core_enc_block_n276) );
  XOR2X1 aes_core_enc_block_U520 ( .A(aes_core_enc_block_n989), .B(
        aes_core_enc_block_n990), .Y(aes_core_enc_block_n988) );
  XOR2X1 aes_core_enc_block_U519 ( .A(aes_core_enc_block_n509), .B(
        aes_core_enc_block_n510), .Y(aes_core_enc_block_n508) );
  XOR2X1 aes_core_enc_block_U518 ( .A(aes_core_enc_block_n750), .B(
        aes_core_enc_block_n751), .Y(aes_core_enc_block_n749) );
  XOR2X1 aes_core_enc_block_U517 ( .A(aes_core_enc_block_n979), .B(
        aes_core_enc_block_n980), .Y(aes_core_enc_block_n978) );
  XOR2X1 aes_core_enc_block_U516 ( .A(aes_core_enc_block_n971), .B(
        aes_core_enc_block_n972), .Y(aes_core_enc_block_n970) );
  XOR2X1 aes_core_enc_block_U515 ( .A(aes_core_enc_block_n732), .B(
        aes_core_enc_block_n733), .Y(aes_core_enc_block_n731) );
  XOR2X1 aes_core_enc_block_U514 ( .A(aes_core_enc_block_n259), .B(
        aes_core_enc_block_n260), .Y(aes_core_enc_block_n258) );
  XOR2X1 aes_core_enc_block_U513 ( .A(aes_core_enc_block_n491), .B(
        aes_core_enc_block_n492), .Y(aes_core_enc_block_n490) );
  XOR2X1 aes_core_enc_block_U512 ( .A(aes_core_enc_block_n294), .B(
        aes_core_enc_block_n295), .Y(aes_core_enc_block_n293) );
  XOR2X1 aes_core_enc_block_U511 ( .A(aes_core_enc_block_n1006), .B(
        aes_core_enc_block_n1007), .Y(aes_core_enc_block_n1005) );
  XOR2X1 aes_core_enc_block_U510 ( .A(aes_core_enc_block_n767), .B(
        aes_core_enc_block_n768), .Y(aes_core_enc_block_n766) );
  XOR2X1 aes_core_enc_block_U509 ( .A(aes_core_enc_block_n526), .B(
        aes_core_enc_block_n527), .Y(aes_core_enc_block_n525) );
  XOR2X1 aes_core_enc_block_U508 ( .A(aes_core_enc_block_n741), .B(
        aes_core_enc_block_n776), .Y(aes_core_enc_block_n775) );
  XOR2X1 aes_core_enc_block_U507 ( .A(aes_core_enc_block_n268), .B(
        aes_core_enc_block_n303), .Y(aes_core_enc_block_n302) );
  XOR2X1 aes_core_enc_block_U506 ( .A(aes_core_enc_block_n980), .B(
        aes_core_enc_block_n1015), .Y(aes_core_enc_block_n1014) );
  XOR2X1 aes_core_enc_block_U505 ( .A(aes_core_enc_block_n500), .B(
        aes_core_enc_block_n535), .Y(aes_core_enc_block_n534) );
  NAND2X1 aes_core_enc_block_U504 ( .A(aes_core_enc_block_n1195), .B(
        aes_core_enc_block_n172), .Y(aes_core_enc_block_n1206) );
  OAI2BB2X1 aes_core_enc_block_U503 ( .B0(aes_core_enc_block_n1204), .B1(
        aes_core_enc_block_n184), .A0N(aes_core_enc_block_n184), .A1N(
        aes_core_enc_block_n1200), .Y(aes_core_enc_block_n1341) );
  AOI21X1 aes_core_enc_block_U502 ( .A0(aes_core_enc_block_n707), .A1(
        aes_core_enc_block_n176), .B0(aes_core_enc_block_n946), .Y(
        aes_core_enc_block_n1208) );
  OAI22X1 aes_core_enc_block_U501 ( .A0(aes_core_enc_block_n174), .A1(
        aes_core_enc_block_n176), .B0(aes_core_enc_block_n1208), .B1(
        aes_core_enc_block_n177), .Y(aes_core_enc_block_n1345) );
  NAND2X1 aes_core_enc_block_U500 ( .A(aes_core_enc_block_n1203), .B(
        aes_core_enc_block_n1196), .Y(aes_core_enc_block_n1205) );
  NOR2X1 aes_core_enc_block_U499 ( .A(aes_core_enc_block_n177), .B(
        aes_core_enc_block_n1195), .Y(aes_core_enc_block_n1209) );
  OAI211X1 aes_core_enc_block_U498 ( .A0(aes_core_enc_block_n172), .A1(
        aes_core_enc_block_n181), .B0(aes_core_enc_block_n1196), .C0(
        aes_core_enc_block_n1206), .Y(aes_core_enc_block_n1343) );
  OAI211X1 aes_core_enc_block_U497 ( .A0(aes_core_enc_block_n172), .A1(
        aes_core_enc_block_n180), .B0(aes_core_enc_block_n1206), .C0(
        aes_core_enc_block_n1193), .Y(aes_core_enc_block_n1344) );
  INVX1 aes_core_enc_block_U496 ( .A(aes_core_enc_block_n1205), .Y(
        aes_core_enc_block_n178) );
  AOI21X1 aes_core_enc_block_U495 ( .A0(aes_core_enc_block_n182), .A1(
        aes_core_enc_block_n177), .B0(aes_core_enc_block_n178), .Y(
        aes_core_enc_block_n1204) );
  INVX1 aes_core_enc_block_U494 ( .A(aes_core_enc_block_n1203), .Y(
        aes_core_enc_block_n177) );
  XNOR2X1 aes_core_enc_block_U493 ( .A(aes_core_round_key[96]), .B(
        aes_core_enc_block_n1423), .Y(aes_core_enc_block_n1190) );
  XOR2X1 aes_core_enc_block_U492 ( .A(aes_core_enc_block_n295), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n1191) );
  XOR2X1 aes_core_enc_block_U491 ( .A(aes_core_enc_block_n1190), .B(
        aes_core_enc_block_n1191), .Y(aes_core_enc_block_n1189) );
  XNOR2X1 aes_core_enc_block_U490 ( .A(aes_core_round_key[42]), .B(
        aes_core_enc_block_n1347), .Y(aes_core_enc_block_n873) );
  XOR2X1 aes_core_enc_block_U489 ( .A(aes_core_enc_block_n751), .B(
        aes_core_enc_block_n767), .Y(aes_core_enc_block_n874) );
  XOR2X1 aes_core_enc_block_U488 ( .A(aes_core_enc_block_n873), .B(
        aes_core_enc_block_n874), .Y(aes_core_enc_block_n872) );
  XNOR2X1 aes_core_enc_block_U487 ( .A(aes_core_round_key[109]), .B(
        aes_core_enc_block_n195), .Y(aes_core_enc_block_n379) );
  XOR2X1 aes_core_enc_block_U486 ( .A(aes_core_enc_block_n252), .B(
        aes_core_enc_block_n269), .Y(aes_core_enc_block_n380) );
  XOR2X1 aes_core_enc_block_U485 ( .A(aes_core_enc_block_n379), .B(
        aes_core_enc_block_n380), .Y(aes_core_enc_block_n378) );
  XNOR2X1 aes_core_enc_block_U484 ( .A(aes_core_round_key[5]), .B(
        aes_core_enc_block_n1404), .Y(aes_core_enc_block_n1147) );
  XNOR2X1 aes_core_enc_block_U483 ( .A(aes_core_enc_block_n1350), .B(
        aes_core_enc_block_n1147), .Y(aes_core_enc_block_n1145) );
  XNOR2X1 aes_core_enc_block_U482 ( .A(aes_core_enc_block_n1389), .B(
        aes_core_enc_block_n964), .Y(aes_core_enc_block_n1146) );
  XOR2X1 aes_core_enc_block_U481 ( .A(aes_core_enc_block_n1145), .B(
        aes_core_enc_block_n1146), .Y(aes_core_enc_block_n1144) );
  XNOR2X1 aes_core_enc_block_U480 ( .A(aes_core_round_key[110]), .B(
        aes_core_enc_block_n240), .Y(aes_core_enc_block_n373) );
  XOR2X1 aes_core_enc_block_U479 ( .A(aes_core_enc_block_n243), .B(
        aes_core_enc_block_n259), .Y(aes_core_enc_block_n374) );
  XOR2X1 aes_core_enc_block_U478 ( .A(aes_core_enc_block_n373), .B(
        aes_core_enc_block_n374), .Y(aes_core_enc_block_n372) );
  XNOR2X1 aes_core_enc_block_U477 ( .A(aes_core_round_key[6]), .B(
        aes_core_enc_block_n1370), .Y(aes_core_enc_block_n1140) );
  XNOR2X1 aes_core_enc_block_U476 ( .A(aes_core_enc_block_n194), .B(
        aes_core_enc_block_n1140), .Y(aes_core_enc_block_n1138) );
  XNOR2X1 aes_core_enc_block_U475 ( .A(aes_core_enc_block_n1379), .B(
        aes_core_enc_block_n955), .Y(aes_core_enc_block_n1139) );
  XOR2X1 aes_core_enc_block_U474 ( .A(aes_core_enc_block_n1138), .B(
        aes_core_enc_block_n1139), .Y(aes_core_enc_block_n1137) );
  XNOR2X1 aes_core_enc_block_U473 ( .A(aes_core_round_key[111]), .B(
        aes_core_enc_block_n1417), .Y(aes_core_enc_block_n367) );
  XOR2X1 aes_core_enc_block_U472 ( .A(aes_core_enc_block_n251), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n368) );
  XOR2X1 aes_core_enc_block_U471 ( .A(aes_core_enc_block_n367), .B(
        aes_core_enc_block_n368), .Y(aes_core_enc_block_n366) );
  XNOR2X1 aes_core_enc_block_U470 ( .A(aes_core_round_key[39]), .B(
        aes_core_enc_block_n1358), .Y(aes_core_enc_block_n894) );
  XNOR2X1 aes_core_enc_block_U469 ( .A(aes_core_enc_block_n1394), .B(
        aes_core_enc_block_n894), .Y(aes_core_enc_block_n892) );
  XNOR2X1 aes_core_enc_block_U468 ( .A(aes_core_enc_block_n1393), .B(
        aes_core_enc_block_n717), .Y(aes_core_enc_block_n893) );
  XOR2X1 aes_core_enc_block_U467 ( .A(aes_core_enc_block_n892), .B(
        aes_core_enc_block_n893), .Y(aes_core_enc_block_n891) );
  XNOR2X1 aes_core_enc_block_U466 ( .A(aes_core_round_key[66]), .B(
        aes_core_enc_block_n1207), .Y(aes_core_enc_block_n690) );
  XNOR2X1 aes_core_enc_block_U465 ( .A(aes_core_enc_block_n1432), .B(
        aes_core_enc_block_n690), .Y(aes_core_enc_block_n688) );
  XNOR2X1 aes_core_enc_block_U464 ( .A(aes_core_enc_block_n1458), .B(
        aes_core_enc_block_n510), .Y(aes_core_enc_block_n689) );
  XOR2X1 aes_core_enc_block_U463 ( .A(aes_core_enc_block_n688), .B(
        aes_core_enc_block_n689), .Y(aes_core_enc_block_n687) );
  XNOR2X1 aes_core_enc_block_U462 ( .A(aes_core_round_key[43]), .B(
        aes_core_enc_block_n1376), .Y(aes_core_enc_block_n868) );
  XOR2X1 aes_core_enc_block_U461 ( .A(aes_core_enc_block_n740), .B(
        aes_core_enc_block_n868), .Y(aes_core_enc_block_n866) );
  XOR2X1 aes_core_enc_block_U460 ( .A(aes_core_enc_block_n759), .B(
        aes_core_enc_block_n860), .Y(aes_core_enc_block_n867) );
  XOR2X1 aes_core_enc_block_U459 ( .A(aes_core_enc_block_n866), .B(
        aes_core_enc_block_n867), .Y(aes_core_enc_block_n865) );
  XNOR2X1 aes_core_enc_block_U458 ( .A(aes_core_round_key[108]), .B(
        aes_core_enc_block_n192), .Y(aes_core_enc_block_n388) );
  XOR2X1 aes_core_enc_block_U457 ( .A(aes_core_enc_block_n260), .B(
        aes_core_enc_block_n388), .Y(aes_core_enc_block_n385) );
  XOR2X1 aes_core_enc_block_U456 ( .A(aes_core_enc_block_n277), .B(
        aes_core_enc_block_n387), .Y(aes_core_enc_block_n386) );
  XOR2X1 aes_core_enc_block_U455 ( .A(aes_core_enc_block_n385), .B(
        aes_core_enc_block_n386), .Y(aes_core_enc_block_n384) );
  XNOR2X1 aes_core_enc_block_U454 ( .A(aes_core_round_key[12]), .B(
        aes_core_enc_block_n1350), .Y(aes_core_enc_block_n1100) );
  XOR2X1 aes_core_enc_block_U453 ( .A(aes_core_enc_block_n972), .B(
        aes_core_enc_block_n1100), .Y(aes_core_enc_block_n1097) );
  XOR2X1 aes_core_enc_block_U452 ( .A(aes_core_enc_block_n989), .B(
        aes_core_enc_block_n1099), .Y(aes_core_enc_block_n1098) );
  XOR2X1 aes_core_enc_block_U451 ( .A(aes_core_enc_block_n1097), .B(
        aes_core_enc_block_n1098), .Y(aes_core_enc_block_n1096) );
  XNOR2X1 aes_core_enc_block_U450 ( .A(aes_core_round_key[45]), .B(
        aes_core_enc_block_n1355), .Y(aes_core_enc_block_n852) );
  XOR2X1 aes_core_enc_block_U449 ( .A(aes_core_enc_block_n725), .B(
        aes_core_enc_block_n742), .Y(aes_core_enc_block_n853) );
  XOR2X1 aes_core_enc_block_U448 ( .A(aes_core_enc_block_n852), .B(
        aes_core_enc_block_n853), .Y(aes_core_enc_block_n851) );
  XNOR2X1 aes_core_enc_block_U447 ( .A(aes_core_round_key[101]), .B(
        aes_core_enc_block_n192), .Y(aes_core_enc_block_n435) );
  XNOR2X1 aes_core_enc_block_U446 ( .A(aes_core_enc_block_n1353), .B(
        aes_core_enc_block_n435), .Y(aes_core_enc_block_n433) );
  XNOR2X1 aes_core_enc_block_U445 ( .A(aes_core_enc_block_n1387), .B(
        aes_core_enc_block_n252), .Y(aes_core_enc_block_n434) );
  XOR2X1 aes_core_enc_block_U444 ( .A(aes_core_enc_block_n433), .B(
        aes_core_enc_block_n434), .Y(aes_core_enc_block_n432) );
  XNOR2X1 aes_core_enc_block_U443 ( .A(aes_core_round_key[69]), .B(
        aes_core_enc_block_n1402), .Y(aes_core_enc_block_n667) );
  XNOR2X1 aes_core_enc_block_U442 ( .A(aes_core_enc_block_n1369), .B(
        aes_core_enc_block_n667), .Y(aes_core_enc_block_n665) );
  XNOR2X1 aes_core_enc_block_U441 ( .A(aes_core_enc_block_n1367), .B(
        aes_core_enc_block_n484), .Y(aes_core_enc_block_n666) );
  XOR2X1 aes_core_enc_block_U440 ( .A(aes_core_enc_block_n665), .B(
        aes_core_enc_block_n666), .Y(aes_core_enc_block_n664) );
  XNOR2X1 aes_core_enc_block_U439 ( .A(aes_core_round_key[46]), .B(
        aes_core_enc_block_n1358), .Y(aes_core_enc_block_n846) );
  XOR2X1 aes_core_enc_block_U438 ( .A(aes_core_enc_block_n716), .B(
        aes_core_enc_block_n732), .Y(aes_core_enc_block_n847) );
  XOR2X1 aes_core_enc_block_U437 ( .A(aes_core_enc_block_n846), .B(
        aes_core_enc_block_n847), .Y(aes_core_enc_block_n845) );
  XNOR2X1 aes_core_enc_block_U436 ( .A(aes_core_round_key[102]), .B(
        aes_core_enc_block_n195), .Y(aes_core_enc_block_n428) );
  XNOR2X1 aes_core_enc_block_U435 ( .A(aes_core_enc_block_n1356), .B(
        aes_core_enc_block_n428), .Y(aes_core_enc_block_n426) );
  XNOR2X1 aes_core_enc_block_U434 ( .A(aes_core_enc_block_n1408), .B(
        aes_core_enc_block_n243), .Y(aes_core_enc_block_n427) );
  XOR2X1 aes_core_enc_block_U433 ( .A(aes_core_enc_block_n426), .B(
        aes_core_enc_block_n427), .Y(aes_core_enc_block_n425) );
  XNOR2X1 aes_core_enc_block_U432 ( .A(aes_core_round_key[70]), .B(
        aes_core_enc_block_n1403), .Y(aes_core_enc_block_n660) );
  XNOR2X1 aes_core_enc_block_U431 ( .A(aes_core_enc_block_n1381), .B(
        aes_core_enc_block_n660), .Y(aes_core_enc_block_n658) );
  XNOR2X1 aes_core_enc_block_U430 ( .A(aes_core_enc_block_n1354), .B(
        aes_core_enc_block_n475), .Y(aes_core_enc_block_n659) );
  XOR2X1 aes_core_enc_block_U429 ( .A(aes_core_enc_block_n658), .B(
        aes_core_enc_block_n659), .Y(aes_core_enc_block_n657) );
  XNOR2X1 aes_core_enc_block_U428 ( .A(aes_core_round_key[47]), .B(
        aes_core_enc_block_n1419), .Y(aes_core_enc_block_n840) );
  XOR2X1 aes_core_enc_block_U427 ( .A(aes_core_enc_block_n724), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n841) );
  XOR2X1 aes_core_enc_block_U426 ( .A(aes_core_enc_block_n840), .B(
        aes_core_enc_block_n841), .Y(aes_core_enc_block_n839) );
  XNOR2X1 aes_core_enc_block_U425 ( .A(aes_core_round_key[103]), .B(
        aes_core_enc_block_n240), .Y(aes_core_enc_block_n421) );
  XNOR2X1 aes_core_enc_block_U424 ( .A(aes_core_enc_block_n1420), .B(
        aes_core_enc_block_n421), .Y(aes_core_enc_block_n419) );
  XNOR2X1 aes_core_enc_block_U423 ( .A(aes_core_enc_block_n1409), .B(
        aes_core_enc_block_n244), .Y(aes_core_enc_block_n420) );
  XOR2X1 aes_core_enc_block_U422 ( .A(aes_core_enc_block_n419), .B(
        aes_core_enc_block_n420), .Y(aes_core_enc_block_n418) );
  XNOR2X1 aes_core_enc_block_U421 ( .A(aes_core_round_key[64]), .B(
        aes_core_enc_block_n1428), .Y(aes_core_enc_block_n703) );
  XOR2X1 aes_core_enc_block_U420 ( .A(aes_core_enc_block_n527), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n704) );
  XOR2X1 aes_core_enc_block_U419 ( .A(aes_core_enc_block_n703), .B(
        aes_core_enc_block_n704), .Y(aes_core_enc_block_n702) );
  XNOR2X1 aes_core_enc_block_U418 ( .A(aes_core_round_key[106]), .B(
        aes_core_enc_block_n1457), .Y(aes_core_enc_block_n400) );
  XOR2X1 aes_core_enc_block_U417 ( .A(aes_core_enc_block_n278), .B(
        aes_core_enc_block_n294), .Y(aes_core_enc_block_n401) );
  XOR2X1 aes_core_enc_block_U416 ( .A(aes_core_enc_block_n400), .B(
        aes_core_enc_block_n401), .Y(aes_core_enc_block_n399) );
  XNOR2X1 aes_core_enc_block_U415 ( .A(aes_core_round_key[76]), .B(
        aes_core_enc_block_n1367), .Y(aes_core_enc_block_n620) );
  XOR2X1 aes_core_enc_block_U414 ( .A(aes_core_enc_block_n492), .B(
        aes_core_enc_block_n620), .Y(aes_core_enc_block_n617) );
  XOR2X1 aes_core_enc_block_U413 ( .A(aes_core_enc_block_n509), .B(
        aes_core_enc_block_n619), .Y(aes_core_enc_block_n618) );
  XOR2X1 aes_core_enc_block_U412 ( .A(aes_core_enc_block_n617), .B(
        aes_core_enc_block_n618), .Y(aes_core_enc_block_n616) );
  XNOR2X1 aes_core_enc_block_U411 ( .A(aes_core_round_key[13]), .B(
        aes_core_enc_block_n194), .Y(aes_core_enc_block_n1091) );
  XOR2X1 aes_core_enc_block_U410 ( .A(aes_core_enc_block_n964), .B(
        aes_core_enc_block_n981), .Y(aes_core_enc_block_n1092) );
  XOR2X1 aes_core_enc_block_U409 ( .A(aes_core_enc_block_n1091), .B(
        aes_core_enc_block_n1092), .Y(aes_core_enc_block_n1090) );
  XNOR2X1 aes_core_enc_block_U408 ( .A(aes_core_round_key[78]), .B(
        aes_core_enc_block_n1357), .Y(aes_core_enc_block_n605) );
  XOR2X1 aes_core_enc_block_U407 ( .A(aes_core_enc_block_n475), .B(
        aes_core_enc_block_n491), .Y(aes_core_enc_block_n606) );
  XOR2X1 aes_core_enc_block_U406 ( .A(aes_core_enc_block_n605), .B(
        aes_core_enc_block_n606), .Y(aes_core_enc_block_n604) );
  XNOR2X1 aes_core_enc_block_U405 ( .A(aes_core_round_key[15]), .B(
        aes_core_enc_block_n1418), .Y(aes_core_enc_block_n1079) );
  XOR2X1 aes_core_enc_block_U404 ( .A(aes_core_enc_block_n963), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1080) );
  XOR2X1 aes_core_enc_block_U403 ( .A(aes_core_enc_block_n1079), .B(
        aes_core_enc_block_n1080), .Y(aes_core_enc_block_n1078) );
  XNOR2X1 aes_core_enc_block_U402 ( .A(aes_core_round_key[74]), .B(
        aes_core_enc_block_n1398), .Y(aes_core_enc_block_n632) );
  XOR2X1 aes_core_enc_block_U401 ( .A(aes_core_enc_block_n510), .B(
        aes_core_enc_block_n526), .Y(aes_core_enc_block_n633) );
  XOR2X1 aes_core_enc_block_U400 ( .A(aes_core_enc_block_n632), .B(
        aes_core_enc_block_n633), .Y(aes_core_enc_block_n631) );
  XNOR2X1 aes_core_enc_block_U399 ( .A(aes_core_round_key[11]), .B(
        aes_core_enc_block_n191), .Y(aes_core_enc_block_n1107) );
  XOR2X1 aes_core_enc_block_U398 ( .A(aes_core_enc_block_n979), .B(
        aes_core_enc_block_n1107), .Y(aes_core_enc_block_n1105) );
  XOR2X1 aes_core_enc_block_U397 ( .A(aes_core_enc_block_n998), .B(
        aes_core_enc_block_n1099), .Y(aes_core_enc_block_n1106) );
  XOR2X1 aes_core_enc_block_U396 ( .A(aes_core_enc_block_n1105), .B(
        aes_core_enc_block_n1106), .Y(aes_core_enc_block_n1104) );
  XNOR2X1 aes_core_enc_block_U395 ( .A(aes_core_round_key[44]), .B(
        aes_core_enc_block_n1352), .Y(aes_core_enc_block_n861) );
  XOR2X1 aes_core_enc_block_U394 ( .A(aes_core_enc_block_n733), .B(
        aes_core_enc_block_n861), .Y(aes_core_enc_block_n858) );
  XOR2X1 aes_core_enc_block_U393 ( .A(aes_core_enc_block_n750), .B(
        aes_core_enc_block_n860), .Y(aes_core_enc_block_n859) );
  XOR2X1 aes_core_enc_block_U392 ( .A(aes_core_enc_block_n858), .B(
        aes_core_enc_block_n859), .Y(aes_core_enc_block_n857) );
  XNOR2X1 aes_core_enc_block_U391 ( .A(aes_core_round_key[117]), .B(
        aes_core_enc_block_n1366), .Y(aes_core_enc_block_n325) );
  XNOR2X1 aes_core_enc_block_U390 ( .A(aes_core_enc_block_n1377), .B(
        aes_core_enc_block_n325), .Y(aes_core_enc_block_n323) );
  XNOR2X1 aes_core_enc_block_U389 ( .A(aes_core_enc_block_n1408), .B(
        aes_core_enc_block_n259), .Y(aes_core_enc_block_n324) );
  XOR2X1 aes_core_enc_block_U388 ( .A(aes_core_enc_block_n323), .B(
        aes_core_enc_block_n324), .Y(aes_core_enc_block_n322) );
  XNOR2X1 aes_core_enc_block_U387 ( .A(aes_core_round_key[14]), .B(
        aes_core_enc_block_n232), .Y(aes_core_enc_block_n1085) );
  XOR2X1 aes_core_enc_block_U386 ( .A(aes_core_enc_block_n955), .B(
        aes_core_enc_block_n971), .Y(aes_core_enc_block_n1086) );
  XOR2X1 aes_core_enc_block_U385 ( .A(aes_core_enc_block_n1085), .B(
        aes_core_enc_block_n1086), .Y(aes_core_enc_block_n1084) );
  XNOR2X1 aes_core_enc_block_U384 ( .A(aes_core_round_key[79]), .B(
        aes_core_enc_block_n1416), .Y(aes_core_enc_block_n599) );
  XOR2X1 aes_core_enc_block_U383 ( .A(aes_core_enc_block_n483), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n600) );
  XOR2X1 aes_core_enc_block_U382 ( .A(aes_core_enc_block_n599), .B(
        aes_core_enc_block_n600), .Y(aes_core_enc_block_n598) );
  XNOR2X1 aes_core_enc_block_U381 ( .A(aes_core_round_key[7]), .B(
        aes_core_enc_block_n232), .Y(aes_core_enc_block_n1133) );
  XNOR2X1 aes_core_enc_block_U380 ( .A(aes_core_enc_block_n1383), .B(
        aes_core_enc_block_n1133), .Y(aes_core_enc_block_n1131) );
  XNOR2X1 aes_core_enc_block_U379 ( .A(aes_core_enc_block_n1380), .B(
        aes_core_enc_block_n956), .Y(aes_core_enc_block_n1132) );
  XOR2X1 aes_core_enc_block_U378 ( .A(aes_core_enc_block_n1131), .B(
        aes_core_enc_block_n1132), .Y(aes_core_enc_block_n1130) );
  XNOR2X1 aes_core_enc_block_U377 ( .A(aes_core_round_key[98]), .B(
        aes_core_enc_block_n189), .Y(aes_core_enc_block_n458) );
  XNOR2X1 aes_core_enc_block_U376 ( .A(aes_core_enc_block_n1397), .B(
        aes_core_enc_block_n458), .Y(aes_core_enc_block_n456) );
  XNOR2X1 aes_core_enc_block_U375 ( .A(aes_core_enc_block_n1434), .B(
        aes_core_enc_block_n278), .Y(aes_core_enc_block_n457) );
  XOR2X1 aes_core_enc_block_U374 ( .A(aes_core_enc_block_n456), .B(
        aes_core_enc_block_n457), .Y(aes_core_enc_block_n455) );
  XNOR2X1 aes_core_enc_block_U373 ( .A(aes_core_round_key[75]), .B(
        aes_core_enc_block_n1385), .Y(aes_core_enc_block_n627) );
  XOR2X1 aes_core_enc_block_U372 ( .A(aes_core_enc_block_n499), .B(
        aes_core_enc_block_n627), .Y(aes_core_enc_block_n625) );
  XOR2X1 aes_core_enc_block_U371 ( .A(aes_core_enc_block_n518), .B(
        aes_core_enc_block_n619), .Y(aes_core_enc_block_n626) );
  XOR2X1 aes_core_enc_block_U370 ( .A(aes_core_enc_block_n625), .B(
        aes_core_enc_block_n626), .Y(aes_core_enc_block_n624) );
  XNOR2X1 aes_core_enc_block_U369 ( .A(aes_core_round_key[77]), .B(
        aes_core_enc_block_n1354), .Y(aes_core_enc_block_n611) );
  XOR2X1 aes_core_enc_block_U368 ( .A(aes_core_enc_block_n484), .B(
        aes_core_enc_block_n501), .Y(aes_core_enc_block_n612) );
  XOR2X1 aes_core_enc_block_U367 ( .A(aes_core_enc_block_n611), .B(
        aes_core_enc_block_n612), .Y(aes_core_enc_block_n610) );
  XNOR2X1 aes_core_enc_block_U366 ( .A(aes_core_round_key[21]), .B(
        aes_core_enc_block_n1368), .Y(aes_core_enc_block_n1037) );
  XNOR2X1 aes_core_enc_block_U365 ( .A(aes_core_enc_block_n1379), .B(
        aes_core_enc_block_n1037), .Y(aes_core_enc_block_n1035) );
  XNOR2X1 aes_core_enc_block_U364 ( .A(aes_core_enc_block_n1388), .B(
        aes_core_enc_block_n971), .Y(aes_core_enc_block_n1036) );
  XOR2X1 aes_core_enc_block_U363 ( .A(aes_core_enc_block_n1035), .B(
        aes_core_enc_block_n1036), .Y(aes_core_enc_block_n1034) );
  XNOR2X1 aes_core_enc_block_U362 ( .A(aes_core_round_key[53]), .B(
        aes_core_enc_block_n1392), .Y(aes_core_enc_block_n798) );
  XNOR2X1 aes_core_enc_block_U361 ( .A(aes_core_enc_block_n1390), .B(
        aes_core_enc_block_n798), .Y(aes_core_enc_block_n796) );
  XNOR2X1 aes_core_enc_block_U360 ( .A(aes_core_enc_block_n1349), .B(
        aes_core_enc_block_n732), .Y(aes_core_enc_block_n797) );
  XOR2X1 aes_core_enc_block_U359 ( .A(aes_core_enc_block_n796), .B(
        aes_core_enc_block_n797), .Y(aes_core_enc_block_n795) );
  XNOR2X1 aes_core_enc_block_U358 ( .A(aes_core_round_key[85]), .B(
        aes_core_enc_block_n1403), .Y(aes_core_enc_block_n557) );
  XNOR2X1 aes_core_enc_block_U357 ( .A(aes_core_enc_block_n1401), .B(
        aes_core_enc_block_n557), .Y(aes_core_enc_block_n555) );
  XNOR2X1 aes_core_enc_block_U356 ( .A(aes_core_enc_block_n1351), .B(
        aes_core_enc_block_n491), .Y(aes_core_enc_block_n556) );
  XOR2X1 aes_core_enc_block_U355 ( .A(aes_core_enc_block_n555), .B(
        aes_core_enc_block_n556), .Y(aes_core_enc_block_n554) );
  XNOR2X1 aes_core_enc_block_U354 ( .A(aes_core_round_key[118]), .B(
        aes_core_enc_block_n1407), .Y(aes_core_enc_block_n318) );
  XNOR2X1 aes_core_enc_block_U353 ( .A(aes_core_enc_block_n1353), .B(
        aes_core_enc_block_n318), .Y(aes_core_enc_block_n316) );
  XNOR2X1 aes_core_enc_block_U352 ( .A(aes_core_enc_block_n1409), .B(
        aes_core_enc_block_n251), .Y(aes_core_enc_block_n317) );
  XOR2X1 aes_core_enc_block_U351 ( .A(aes_core_enc_block_n316), .B(
        aes_core_enc_block_n317), .Y(aes_core_enc_block_n315) );
  XNOR2X1 aes_core_enc_block_U350 ( .A(aes_core_round_key[22]), .B(
        aes_core_enc_block_n1404), .Y(aes_core_enc_block_n1030) );
  XNOR2X1 aes_core_enc_block_U349 ( .A(aes_core_enc_block_n1380), .B(
        aes_core_enc_block_n1030), .Y(aes_core_enc_block_n1028) );
  XNOR2X1 aes_core_enc_block_U348 ( .A(aes_core_enc_block_n1378), .B(
        aes_core_enc_block_n963), .Y(aes_core_enc_block_n1029) );
  XOR2X1 aes_core_enc_block_U347 ( .A(aes_core_enc_block_n1028), .B(
        aes_core_enc_block_n1029), .Y(aes_core_enc_block_n1027) );
  XNOR2X1 aes_core_enc_block_U346 ( .A(aes_core_round_key[54]), .B(
        aes_core_enc_block_n1393), .Y(aes_core_enc_block_n791) );
  XNOR2X1 aes_core_enc_block_U345 ( .A(aes_core_enc_block_n1405), .B(
        aes_core_enc_block_n791), .Y(aes_core_enc_block_n789) );
  XNOR2X1 aes_core_enc_block_U344 ( .A(aes_core_enc_block_n193), .B(
        aes_core_enc_block_n724), .Y(aes_core_enc_block_n790) );
  XOR2X1 aes_core_enc_block_U343 ( .A(aes_core_enc_block_n789), .B(
        aes_core_enc_block_n790), .Y(aes_core_enc_block_n788) );
  XNOR2X1 aes_core_enc_block_U342 ( .A(aes_core_round_key[86]), .B(
        aes_core_enc_block_n1413), .Y(aes_core_enc_block_n550) );
  XNOR2X1 aes_core_enc_block_U341 ( .A(aes_core_enc_block_n1406), .B(
        aes_core_enc_block_n550), .Y(aes_core_enc_block_n548) );
  XNOR2X1 aes_core_enc_block_U340 ( .A(aes_core_enc_block_n1369), .B(
        aes_core_enc_block_n483), .Y(aes_core_enc_block_n549) );
  XOR2X1 aes_core_enc_block_U339 ( .A(aes_core_enc_block_n548), .B(
        aes_core_enc_block_n549), .Y(aes_core_enc_block_n547) );
  XNOR2X1 aes_core_enc_block_U338 ( .A(aes_core_round_key[71]), .B(
        aes_core_enc_block_n1361), .Y(aes_core_enc_block_n653) );
  XNOR2X1 aes_core_enc_block_U337 ( .A(aes_core_enc_block_n1413), .B(
        aes_core_enc_block_n653), .Y(aes_core_enc_block_n651) );
  XNOR2X1 aes_core_enc_block_U336 ( .A(aes_core_enc_block_n1357), .B(
        aes_core_enc_block_n476), .Y(aes_core_enc_block_n652) );
  XOR2X1 aes_core_enc_block_U335 ( .A(aes_core_enc_block_n651), .B(
        aes_core_enc_block_n652), .Y(aes_core_enc_block_n650) );
  XNOR2X1 aes_core_enc_block_U334 ( .A(aes_core_round_key[55]), .B(
        aes_core_enc_block_n1411), .Y(aes_core_enc_block_n784) );
  XNOR2X1 aes_core_enc_block_U333 ( .A(aes_core_enc_block_n467), .B(
        aes_core_enc_block_n784), .Y(aes_core_enc_block_n781) );
  XNOR2X1 aes_core_enc_block_U332 ( .A(aes_core_enc_block_n196), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n782) );
  XOR2X1 aes_core_enc_block_U331 ( .A(aes_core_enc_block_n781), .B(
        aes_core_enc_block_n782), .Y(aes_core_enc_block_n780) );
  XNOR2X1 aes_core_enc_block_U330 ( .A(aes_core_round_key[87]), .B(
        aes_core_enc_block_n1412), .Y(aes_core_enc_block_n543) );
  XNOR2X1 aes_core_enc_block_U329 ( .A(aes_core_enc_block_n1371), .B(
        aes_core_enc_block_n543), .Y(aes_core_enc_block_n540) );
  XNOR2X1 aes_core_enc_block_U328 ( .A(aes_core_enc_block_n1381), .B(
        aes_core_enc_block_n542), .Y(aes_core_enc_block_n541) );
  XOR2X1 aes_core_enc_block_U327 ( .A(aes_core_enc_block_n540), .B(
        aes_core_enc_block_n541), .Y(aes_core_enc_block_n539) );
  XNOR2X1 aes_core_enc_block_U326 ( .A(aes_core_round_key[119]), .B(
        aes_core_enc_block_n1414), .Y(aes_core_enc_block_n311) );
  XNOR2X1 aes_core_enc_block_U325 ( .A(aes_core_enc_block_n1359), .B(
        aes_core_enc_block_n311), .Y(aes_core_enc_block_n308) );
  XNOR2X1 aes_core_enc_block_U324 ( .A(aes_core_enc_block_n1356), .B(
        aes_core_enc_block_n310), .Y(aes_core_enc_block_n309) );
  XOR2X1 aes_core_enc_block_U323 ( .A(aes_core_enc_block_n308), .B(
        aes_core_enc_block_n309), .Y(aes_core_enc_block_n307) );
  XNOR2X1 aes_core_enc_block_U322 ( .A(aes_core_round_key[23]), .B(
        aes_core_enc_block_n1382), .Y(aes_core_enc_block_n1023) );
  XNOR2X1 aes_core_enc_block_U321 ( .A(aes_core_enc_block_n1370), .B(
        aes_core_enc_block_n1023), .Y(aes_core_enc_block_n1020) );
  XNOR2X1 aes_core_enc_block_U320 ( .A(aes_core_enc_block_n1410), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1021) );
  XOR2X1 aes_core_enc_block_U319 ( .A(aes_core_enc_block_n1020), .B(
        aes_core_enc_block_n1021), .Y(aes_core_enc_block_n1019) );
  XNOR2X1 aes_core_enc_block_U318 ( .A(aes_core_round_key[104]), .B(
        aes_core_enc_block_n947), .Y(aes_core_enc_block_n413) );
  XOR2X1 aes_core_enc_block_U317 ( .A(aes_core_enc_block_n295), .B(
        aes_core_enc_block_n387), .Y(aes_core_enc_block_n414) );
  XOR2X1 aes_core_enc_block_U316 ( .A(aes_core_enc_block_n413), .B(
        aes_core_enc_block_n414), .Y(aes_core_enc_block_n412) );
  XNOR2X1 aes_core_enc_block_U315 ( .A(aes_core_round_key[105]), .B(
        aes_core_enc_block_n1397), .Y(aes_core_enc_block_n408) );
  XOR2X1 aes_core_enc_block_U314 ( .A(aes_core_enc_block_n287), .B(
        aes_core_enc_block_n408), .Y(aes_core_enc_block_n406) );
  XOR2X1 aes_core_enc_block_U313 ( .A(aes_core_enc_block_n303), .B(
        aes_core_enc_block_n387), .Y(aes_core_enc_block_n407) );
  XOR2X1 aes_core_enc_block_U312 ( .A(aes_core_enc_block_n406), .B(
        aes_core_enc_block_n407), .Y(aes_core_enc_block_n405) );
  XNOR2X1 aes_core_enc_block_U311 ( .A(aes_core_round_key[50]), .B(
        aes_core_enc_block_n1441), .Y(aes_core_enc_block_n821) );
  XNOR2X1 aes_core_enc_block_U310 ( .A(aes_core_enc_block_n1439), .B(
        aes_core_enc_block_n821), .Y(aes_core_enc_block_n819) );
  XNOR2X1 aes_core_enc_block_U309 ( .A(aes_core_enc_block_n1436), .B(
        aes_core_enc_block_n759), .Y(aes_core_enc_block_n820) );
  XOR2X1 aes_core_enc_block_U308 ( .A(aes_core_enc_block_n819), .B(
        aes_core_enc_block_n820), .Y(aes_core_enc_block_n818) );
  XNOR2X1 aes_core_enc_block_U307 ( .A(aes_core_round_key[82]), .B(
        aes_core_enc_block_n1373), .Y(aes_core_enc_block_n580) );
  XNOR2X1 aes_core_enc_block_U306 ( .A(aes_core_enc_block_n1443), .B(
        aes_core_enc_block_n580), .Y(aes_core_enc_block_n578) );
  XNOR2X1 aes_core_enc_block_U305 ( .A(aes_core_enc_block_n1431), .B(
        aes_core_enc_block_n518), .Y(aes_core_enc_block_n579) );
  XOR2X1 aes_core_enc_block_U304 ( .A(aes_core_enc_block_n578), .B(
        aes_core_enc_block_n579), .Y(aes_core_enc_block_n577) );
  XNOR2X1 aes_core_enc_block_U303 ( .A(aes_core_round_key[114]), .B(
        aes_core_enc_block_n1433), .Y(aes_core_enc_block_n348) );
  XNOR2X1 aes_core_enc_block_U302 ( .A(aes_core_enc_block_n1363), .B(
        aes_core_enc_block_n348), .Y(aes_core_enc_block_n346) );
  XNOR2X1 aes_core_enc_block_U301 ( .A(aes_core_enc_block_n1445), .B(
        aes_core_enc_block_n286), .Y(aes_core_enc_block_n347) );
  XOR2X1 aes_core_enc_block_U300 ( .A(aes_core_enc_block_n346), .B(
        aes_core_enc_block_n347), .Y(aes_core_enc_block_n345) );
  XNOR2X1 aes_core_enc_block_U299 ( .A(aes_core_round_key[18]), .B(
        aes_core_enc_block_n1437), .Y(aes_core_enc_block_n1060) );
  XNOR2X1 aes_core_enc_block_U298 ( .A(aes_core_enc_block_n1447), .B(
        aes_core_enc_block_n1060), .Y(aes_core_enc_block_n1058) );
  XNOR2X1 aes_core_enc_block_U297 ( .A(aes_core_enc_block_n1435), .B(
        aes_core_enc_block_n998), .Y(aes_core_enc_block_n1059) );
  XOR2X1 aes_core_enc_block_U296 ( .A(aes_core_enc_block_n1058), .B(
        aes_core_enc_block_n1059), .Y(aes_core_enc_block_n1057) );
  XNOR2X1 aes_core_enc_block_U295 ( .A(aes_core_round_key[2]), .B(
        aes_core_enc_block_n1374), .Y(aes_core_enc_block_n1170) );
  XNOR2X1 aes_core_enc_block_U294 ( .A(aes_core_enc_block_n1456), .B(
        aes_core_enc_block_n1170), .Y(aes_core_enc_block_n1168) );
  XNOR2X1 aes_core_enc_block_U293 ( .A(aes_core_enc_block_n1438), .B(
        aes_core_enc_block_n990), .Y(aes_core_enc_block_n1169) );
  XOR2X1 aes_core_enc_block_U292 ( .A(aes_core_enc_block_n1168), .B(
        aes_core_enc_block_n1169), .Y(aes_core_enc_block_n1167) );
  XNOR2X1 aes_core_enc_block_U291 ( .A(aes_core_round_key[10]), .B(
        aes_core_enc_block_n1454), .Y(aes_core_enc_block_n1112) );
  XOR2X1 aes_core_enc_block_U290 ( .A(aes_core_enc_block_n990), .B(
        aes_core_enc_block_n1006), .Y(aes_core_enc_block_n1113) );
  XOR2X1 aes_core_enc_block_U289 ( .A(aes_core_enc_block_n1112), .B(
        aes_core_enc_block_n1113), .Y(aes_core_enc_block_n1111) );
  XNOR2X1 aes_core_enc_block_U288 ( .A(aes_core_round_key[112]), .B(
        aes_core_enc_block_n1421), .Y(aes_core_enc_block_n361) );
  XOR2X1 aes_core_enc_block_U287 ( .A(aes_core_enc_block_n244), .B(
        aes_core_enc_block_n303), .Y(aes_core_enc_block_n362) );
  XOR2X1 aes_core_enc_block_U286 ( .A(aes_core_enc_block_n361), .B(
        aes_core_enc_block_n362), .Y(aes_core_enc_block_n360) );
  XNOR2X1 aes_core_enc_block_U285 ( .A(aes_core_round_key[0]), .B(
        aes_core_enc_block_n1372), .Y(aes_core_enc_block_n1183) );
  XOR2X1 aes_core_enc_block_U284 ( .A(aes_core_enc_block_n1007), .B(
        aes_core_enc_block_n1022), .Y(aes_core_enc_block_n1184) );
  XOR2X1 aes_core_enc_block_U283 ( .A(aes_core_enc_block_n1183), .B(
        aes_core_enc_block_n1184), .Y(aes_core_enc_block_n1182) );
  XNOR2X1 aes_core_enc_block_U282 ( .A(aes_core_round_key[72]), .B(
        aes_core_enc_block_n187), .Y(aes_core_enc_block_n645) );
  XOR2X1 aes_core_enc_block_U281 ( .A(aes_core_enc_block_n527), .B(
        aes_core_enc_block_n619), .Y(aes_core_enc_block_n646) );
  XOR2X1 aes_core_enc_block_U280 ( .A(aes_core_enc_block_n645), .B(
        aes_core_enc_block_n646), .Y(aes_core_enc_block_n644) );
  XNOR2X1 aes_core_enc_block_U279 ( .A(aes_core_round_key[32]), .B(
        aes_core_enc_block_n1422), .Y(aes_core_enc_block_n944) );
  XOR2X1 aes_core_enc_block_U278 ( .A(aes_core_enc_block_n768), .B(
        aes_core_enc_block_n783), .Y(aes_core_enc_block_n945) );
  XOR2X1 aes_core_enc_block_U277 ( .A(aes_core_enc_block_n944), .B(
        aes_core_enc_block_n945), .Y(aes_core_enc_block_n943) );
  XNOR2X1 aes_core_enc_block_U276 ( .A(aes_core_round_key[40]), .B(
        aes_core_enc_block_n1362), .Y(aes_core_enc_block_n886) );
  XOR2X1 aes_core_enc_block_U275 ( .A(aes_core_enc_block_n768), .B(
        aes_core_enc_block_n860), .Y(aes_core_enc_block_n887) );
  XOR2X1 aes_core_enc_block_U274 ( .A(aes_core_enc_block_n886), .B(
        aes_core_enc_block_n887), .Y(aes_core_enc_block_n885) );
  XNOR2X1 aes_core_enc_block_U273 ( .A(aes_core_round_key[16]), .B(
        aes_core_enc_block_n1425), .Y(aes_core_enc_block_n1073) );
  XOR2X1 aes_core_enc_block_U272 ( .A(aes_core_enc_block_n956), .B(
        aes_core_enc_block_n1015), .Y(aes_core_enc_block_n1074) );
  XOR2X1 aes_core_enc_block_U271 ( .A(aes_core_enc_block_n1073), .B(
        aes_core_enc_block_n1074), .Y(aes_core_enc_block_n1072) );
  XNOR2X1 aes_core_enc_block_U270 ( .A(aes_core_round_key[48]), .B(
        aes_core_enc_block_n1395), .Y(aes_core_enc_block_n834) );
  XOR2X1 aes_core_enc_block_U269 ( .A(aes_core_enc_block_n717), .B(
        aes_core_enc_block_n776), .Y(aes_core_enc_block_n835) );
  XOR2X1 aes_core_enc_block_U268 ( .A(aes_core_enc_block_n834), .B(
        aes_core_enc_block_n835), .Y(aes_core_enc_block_n833) );
  XNOR2X1 aes_core_enc_block_U267 ( .A(aes_core_round_key[8]), .B(
        aes_core_enc_block_n1396), .Y(aes_core_enc_block_n1125) );
  XOR2X1 aes_core_enc_block_U266 ( .A(aes_core_enc_block_n1007), .B(
        aes_core_enc_block_n1099), .Y(aes_core_enc_block_n1126) );
  XOR2X1 aes_core_enc_block_U265 ( .A(aes_core_enc_block_n1125), .B(
        aes_core_enc_block_n1126), .Y(aes_core_enc_block_n1124) );
  XNOR2X1 aes_core_enc_block_U264 ( .A(aes_core_round_key[80]), .B(
        aes_core_enc_block_n1429), .Y(aes_core_enc_block_n593) );
  XOR2X1 aes_core_enc_block_U263 ( .A(aes_core_enc_block_n476), .B(
        aes_core_enc_block_n535), .Y(aes_core_enc_block_n594) );
  XOR2X1 aes_core_enc_block_U262 ( .A(aes_core_enc_block_n593), .B(
        aes_core_enc_block_n594), .Y(aes_core_enc_block_n592) );
  XNOR2X1 aes_core_enc_block_U261 ( .A(aes_core_round_key[41]), .B(
        aes_core_enc_block_n188), .Y(aes_core_enc_block_n881) );
  XOR2X1 aes_core_enc_block_U260 ( .A(aes_core_enc_block_n760), .B(
        aes_core_enc_block_n881), .Y(aes_core_enc_block_n879) );
  XOR2X1 aes_core_enc_block_U259 ( .A(aes_core_enc_block_n776), .B(
        aes_core_enc_block_n860), .Y(aes_core_enc_block_n880) );
  XOR2X1 aes_core_enc_block_U258 ( .A(aes_core_enc_block_n879), .B(
        aes_core_enc_block_n880), .Y(aes_core_enc_block_n878) );
  XNOR2X1 aes_core_enc_block_U257 ( .A(aes_core_round_key[9]), .B(
        aes_core_enc_block_n1456), .Y(aes_core_enc_block_n1120) );
  XOR2X1 aes_core_enc_block_U256 ( .A(aes_core_enc_block_n999), .B(
        aes_core_enc_block_n1120), .Y(aes_core_enc_block_n1118) );
  XOR2X1 aes_core_enc_block_U255 ( .A(aes_core_enc_block_n1015), .B(
        aes_core_enc_block_n1099), .Y(aes_core_enc_block_n1119) );
  XOR2X1 aes_core_enc_block_U254 ( .A(aes_core_enc_block_n1118), .B(
        aes_core_enc_block_n1119), .Y(aes_core_enc_block_n1117) );
  XNOR2X1 aes_core_enc_block_U253 ( .A(aes_core_round_key[73]), .B(
        aes_core_enc_block_n1207), .Y(aes_core_enc_block_n640) );
  XOR2X1 aes_core_enc_block_U252 ( .A(aes_core_enc_block_n519), .B(
        aes_core_enc_block_n640), .Y(aes_core_enc_block_n638) );
  XOR2X1 aes_core_enc_block_U251 ( .A(aes_core_enc_block_n535), .B(
        aes_core_enc_block_n619), .Y(aes_core_enc_block_n639) );
  XOR2X1 aes_core_enc_block_U250 ( .A(aes_core_enc_block_n638), .B(
        aes_core_enc_block_n639), .Y(aes_core_enc_block_n637) );
  XNOR2X1 aes_core_enc_block_U249 ( .A(aes_core_round_key[37]), .B(
        aes_core_enc_block_n1352), .Y(aes_core_enc_block_n908) );
  XNOR2X1 aes_core_enc_block_U248 ( .A(aes_core_enc_block_n1391), .B(
        aes_core_enc_block_n908), .Y(aes_core_enc_block_n906) );
  XNOR2X1 aes_core_enc_block_U247 ( .A(aes_core_enc_block_n193), .B(
        aes_core_enc_block_n725), .Y(aes_core_enc_block_n907) );
  XOR2X1 aes_core_enc_block_U246 ( .A(aes_core_enc_block_n906), .B(
        aes_core_enc_block_n907), .Y(aes_core_enc_block_n905) );
  XNOR2X1 aes_core_enc_block_U245 ( .A(aes_core_round_key[38]), .B(
        aes_core_enc_block_n1355), .Y(aes_core_enc_block_n901) );
  XNOR2X1 aes_core_enc_block_U244 ( .A(aes_core_enc_block_n1392), .B(
        aes_core_enc_block_n901), .Y(aes_core_enc_block_n899) );
  XNOR2X1 aes_core_enc_block_U243 ( .A(aes_core_enc_block_n196), .B(
        aes_core_enc_block_n716), .Y(aes_core_enc_block_n900) );
  XOR2X1 aes_core_enc_block_U242 ( .A(aes_core_enc_block_n899), .B(
        aes_core_enc_block_n900), .Y(aes_core_enc_block_n898) );
  XNOR2X1 aes_core_enc_block_U241 ( .A(aes_core_round_key[34]), .B(
        aes_core_enc_block_n188), .Y(aes_core_enc_block_n931) );
  XNOR2X1 aes_core_enc_block_U240 ( .A(aes_core_enc_block_n1440), .B(
        aes_core_enc_block_n931), .Y(aes_core_enc_block_n929) );
  XNOR2X1 aes_core_enc_block_U239 ( .A(aes_core_enc_block_n1364), .B(
        aes_core_enc_block_n751), .Y(aes_core_enc_block_n930) );
  XOR2X1 aes_core_enc_block_U238 ( .A(aes_core_enc_block_n929), .B(
        aes_core_enc_block_n930), .Y(aes_core_enc_block_n928) );
  XNOR2X1 aes_core_enc_block_U237 ( .A(aes_core_round_key[65]), .B(
        aes_core_enc_block_n1373), .Y(aes_core_enc_block_n698) );
  XNOR2X1 aes_core_enc_block_U236 ( .A(aes_core_round_key[35]), .B(
        aes_core_enc_block_n1347), .Y(aes_core_enc_block_n924) );
  XNOR2X1 aes_core_enc_block_U235 ( .A(aes_core_round_key[4]), .B(
        aes_core_enc_block_n1368), .Y(aes_core_enc_block_n1155) );
  XNOR2X1 aes_core_enc_block_U234 ( .A(aes_core_round_key[97]), .B(
        aes_core_enc_block_n1363), .Y(aes_core_enc_block_n466) );
  XNOR2X1 aes_core_enc_block_U233 ( .A(aes_core_round_key[36]), .B(
        aes_core_enc_block_n1376), .Y(aes_core_enc_block_n916) );
  XNOR2X1 aes_core_enc_block_U232 ( .A(aes_core_round_key[68]), .B(
        aes_core_enc_block_n1385), .Y(aes_core_enc_block_n675) );
  XNOR2X1 aes_core_enc_block_U231 ( .A(aes_core_round_key[51]), .B(
        aes_core_enc_block_n1453), .Y(aes_core_enc_block_n814) );
  XNOR2X1 aes_core_enc_block_U230 ( .A(aes_core_round_key[84]), .B(
        aes_core_enc_block_n1402), .Y(aes_core_enc_block_n565) );
  XNOR2X1 aes_core_enc_block_U229 ( .A(aes_core_round_key[100]), .B(
        aes_core_enc_block_n1377), .Y(aes_core_enc_block_n443) );
  XNOR2X1 aes_core_enc_block_U228 ( .A(aes_core_round_key[67]), .B(
        aes_core_enc_block_n1398), .Y(aes_core_enc_block_n683) );
  XNOR2X1 aes_core_enc_block_U227 ( .A(aes_core_round_key[99]), .B(
        aes_core_enc_block_n1348), .Y(aes_core_enc_block_n451) );
  XNOR2X1 aes_core_enc_block_U226 ( .A(aes_core_round_key[83]), .B(
        aes_core_enc_block_n1452), .Y(aes_core_enc_block_n573) );
  XNOR2X1 aes_core_enc_block_U225 ( .A(aes_core_round_key[116]), .B(
        aes_core_enc_block_n1386), .Y(aes_core_enc_block_n333) );
  XNOR2X1 aes_core_enc_block_U224 ( .A(aes_core_round_key[20]), .B(
        aes_core_enc_block_n1399), .Y(aes_core_enc_block_n1045) );
  XNOR2X1 aes_core_enc_block_U223 ( .A(aes_core_round_key[1]), .B(
        aes_core_enc_block_n1437), .Y(aes_core_enc_block_n1178) );
  XNOR2X1 aes_core_enc_block_U222 ( .A(aes_core_round_key[19]), .B(
        aes_core_enc_block_n1374), .Y(aes_core_enc_block_n1053) );
  XNOR2X1 aes_core_enc_block_U221 ( .A(aes_core_round_key[52]), .B(
        aes_core_enc_block_n1391), .Y(aes_core_enc_block_n806) );
  XNOR2X1 aes_core_enc_block_U220 ( .A(aes_core_round_key[49]), .B(
        aes_core_enc_block_n1440), .Y(aes_core_enc_block_n829) );
  XNOR2X1 aes_core_enc_block_U219 ( .A(aes_core_round_key[81]), .B(
        aes_core_enc_block_n1428), .Y(aes_core_enc_block_n588) );
  XNOR2X1 aes_core_enc_block_U218 ( .A(aes_core_round_key[113]), .B(
        aes_core_enc_block_n1430), .Y(aes_core_enc_block_n356) );
  XNOR2X1 aes_core_enc_block_U217 ( .A(aes_core_round_key[17]), .B(
        aes_core_enc_block_n1372), .Y(aes_core_enc_block_n1068) );
  XNOR2X1 aes_core_enc_block_U216 ( .A(aes_core_round_key[115]), .B(
        aes_core_enc_block_n1444), .Y(aes_core_enc_block_n341) );
  XNOR2X1 aes_core_enc_block_U215 ( .A(aes_core_round_key[3]), .B(
        aes_core_enc_block_n1399), .Y(aes_core_enc_block_n1163) );
  XNOR2X1 aes_core_enc_block_U214 ( .A(aes_core_round_key[33]), .B(
        aes_core_enc_block_n1362), .Y(aes_core_enc_block_n939) );
  XNOR2X1 aes_core_enc_block_U213 ( .A(aes_core_round_key[107]), .B(
        aes_core_enc_block_n1455), .Y(aes_core_enc_block_n395) );
  XOR2X1 aes_core_enc_block_U212 ( .A(aes_core_enc_block_n267), .B(
        aes_core_enc_block_n395), .Y(aes_core_enc_block_n393) );
  XOR2X1 aes_core_enc_block_U211 ( .A(aes_core_enc_block_n286), .B(
        aes_core_enc_block_n387), .Y(aes_core_enc_block_n394) );
  XOR2X1 aes_core_enc_block_U210 ( .A(aes_core_enc_block_n393), .B(
        aes_core_enc_block_n394), .Y(aes_core_enc_block_n392) );
  INVX1 aes_core_enc_block_U209 ( .A(aes_core_round_key[124]), .Y(
        aes_core_enc_block_n135) );
  INVX1 aes_core_enc_block_U208 ( .A(aes_core_round_key[28]), .Y(
        aes_core_enc_block_n167) );
  INVX1 aes_core_enc_block_U207 ( .A(aes_core_round_key[60]), .Y(
        aes_core_enc_block_n151) );
  INVX1 aes_core_enc_block_U206 ( .A(aes_core_round_key[92]), .Y(
        aes_core_enc_block_n143) );
  INVX1 aes_core_enc_block_U205 ( .A(aes_core_round_key[89]), .Y(
        aes_core_enc_block_n146) );
  INVX1 aes_core_enc_block_U204 ( .A(aes_core_round_key[121]), .Y(
        aes_core_enc_block_n138) );
  INVX1 aes_core_enc_block_U203 ( .A(aes_core_round_key[25]), .Y(
        aes_core_enc_block_n170) );
  INVX1 aes_core_enc_block_U202 ( .A(aes_core_round_key[57]), .Y(
        aes_core_enc_block_n154) );
  INVX1 aes_core_enc_block_U201 ( .A(aes_core_round_key[123]), .Y(
        aes_core_enc_block_n136) );
  INVX1 aes_core_enc_block_U200 ( .A(aes_core_round_key[27]), .Y(
        aes_core_enc_block_n168) );
  INVX1 aes_core_enc_block_U199 ( .A(aes_core_round_key[91]), .Y(
        aes_core_enc_block_n144) );
  INVX1 aes_core_enc_block_U198 ( .A(aes_core_round_key[59]), .Y(
        aes_core_enc_block_n152) );
  INVX1 aes_core_enc_block_U197 ( .A(aes_core_round_key[95]), .Y(
        aes_core_enc_block_n140) );
  INVX1 aes_core_enc_block_U196 ( .A(aes_core_round_key[29]), .Y(
        aes_core_enc_block_n166) );
  INVX1 aes_core_enc_block_U195 ( .A(aes_core_round_key[30]), .Y(
        aes_core_enc_block_n165) );
  INVX1 aes_core_enc_block_U194 ( .A(aes_core_round_key[31]), .Y(
        aes_core_enc_block_n156) );
  INVX1 aes_core_enc_block_U193 ( .A(aes_core_round_key[61]), .Y(
        aes_core_enc_block_n150) );
  INVX1 aes_core_enc_block_U192 ( .A(aes_core_round_key[62]), .Y(
        aes_core_enc_block_n149) );
  INVX1 aes_core_enc_block_U191 ( .A(aes_core_round_key[63]), .Y(
        aes_core_enc_block_n148) );
  INVX1 aes_core_enc_block_U190 ( .A(aes_core_round_key[56]), .Y(
        aes_core_enc_block_n155) );
  INVX1 aes_core_enc_block_U189 ( .A(aes_core_round_key[93]), .Y(
        aes_core_enc_block_n142) );
  INVX1 aes_core_enc_block_U188 ( .A(aes_core_round_key[125]), .Y(
        aes_core_enc_block_n134) );
  INVX1 aes_core_enc_block_U187 ( .A(aes_core_round_key[126]), .Y(
        aes_core_enc_block_n133) );
  INVX1 aes_core_enc_block_U186 ( .A(aes_core_round_key[94]), .Y(
        aes_core_enc_block_n141) );
  INVX1 aes_core_enc_block_U185 ( .A(aes_core_round_key[127]), .Y(
        aes_core_enc_block_n132) );
  INVX1 aes_core_enc_block_U184 ( .A(aes_core_round_key[120]), .Y(
        aes_core_enc_block_n139) );
  INVX1 aes_core_enc_block_U183 ( .A(aes_core_round_key[24]), .Y(
        aes_core_enc_block_n171) );
  INVX1 aes_core_enc_block_U182 ( .A(aes_core_round_key[88]), .Y(
        aes_core_enc_block_n147) );
  INVX1 aes_core_enc_block_U181 ( .A(aes_core_round_key[58]), .Y(
        aes_core_enc_block_n153) );
  INVX1 aes_core_enc_block_U180 ( .A(aes_core_round_key[90]), .Y(
        aes_core_enc_block_n145) );
  INVX1 aes_core_enc_block_U179 ( .A(aes_core_round_key[122]), .Y(
        aes_core_enc_block_n137) );
  INVX1 aes_core_enc_block_U178 ( .A(aes_core_round_key[26]), .Y(
        aes_core_enc_block_n169) );
  NOR2X1 aes_core_enc_block_U177 ( .A(aes_core_enc_block_n1193), .B(
        aes_core_enc_block_n1192), .Y(aes_core_enc_block_n235) );
  NOR2X1 aes_core_enc_block_U176 ( .A(aes_core_enc_block_n174), .B(
        aes_core_enc_block_n173), .Y(aes_core_enc_block_n1185) );
  NOR2X1 aes_core_enc_block_U175 ( .A(aes_core_enc_block_n181), .B(
        aes_core_enc_block_n180), .Y(aes_core_enc_block_n1194) );
  INVX1 aes_core_enc_block_U174 ( .A(aes_core_enc_block_n1193), .Y(
        aes_core_enc_block_n179) );
  NAND3X1 aes_core_enc_block_U173 ( .A(aes_core_enc_block_n173), .B(
        aes_core_enc_block_n174), .C(aes_core_enc_block_n705), .Y(
        aes_core_enc_block_n197) );
  AOI21X1 aes_core_enc_block_U172 ( .A0(aes_core_enc_block_n184), .A1(
        aes_core_enc_block_n185), .B0(aes_core_enc_block_n186), .Y(
        aes_core_enc_block_n1197) );
  INVX1 aes_core_enc_block_U171 ( .A(aes_core_enc_block_n1209), .Y(
        aes_core_enc_block_n176) );
  INVX1 aes_core_enc_block_U170 ( .A(aes_core_enc_block_n235), .Y(
        aes_core_enc_block_n122) );
  CLKINVX3 aes_core_enc_block_U169 ( .A(aes_core_enc_block_n122), .Y(
        aes_core_enc_block_n117) );
  NAND2X1 aes_core_enc_block_U168 ( .A(aes_core_enc_block_n706), .B(
        aes_core_enc_block_n230), .Y(aes_core_enc_block_n709) );
  NAND2X1 aes_core_enc_block_U167 ( .A(aes_core_enc_block_n1192), .B(
        aes_core_enc_block_n179), .Y(aes_core_enc_block_n239) );
  INVX1 aes_core_enc_block_U166 ( .A(aes_core_new_sboxw[27]), .Y(
        aes_core_enc_block_n162) );
  INVX1 aes_core_enc_block_U165 ( .A(aes_core_new_sboxw[28]), .Y(
        aes_core_enc_block_n158) );
  INVX1 aes_core_enc_block_U164 ( .A(aes_core_new_sboxw[31]), .Y(
        aes_core_enc_block_n159) );
  INVX1 aes_core_enc_block_U163 ( .A(aes_core_enc_block_n1197), .Y(
        aes_core_enc_block_n183) );
  INVX1 aes_core_enc_block_U162 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n88) );
  INVX1 aes_core_enc_block_U161 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n85) );
  INVX1 aes_core_enc_block_U160 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n89) );
  INVX1 aes_core_enc_block_U159 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n90) );
  INVX1 aes_core_enc_block_U158 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n86) );
  INVX1 aes_core_enc_block_U157 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n87) );
  INVX1 aes_core_enc_block_U156 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n91) );
  CLKINVX3 aes_core_enc_block_U155 ( .A(aes_core_enc_block_n122), .Y(
        aes_core_enc_block_n120) );
  CLKINVX3 aes_core_enc_block_U154 ( .A(aes_core_enc_block_n122), .Y(
        aes_core_enc_block_n118) );
  CLKINVX3 aes_core_enc_block_U153 ( .A(aes_core_enc_block_n122), .Y(
        aes_core_enc_block_n119) );
  CLKINVX3 aes_core_enc_block_U152 ( .A(aes_core_enc_block_n122), .Y(
        aes_core_enc_block_n121) );
  INVX1 aes_core_enc_block_U151 ( .A(aes_core_enc_block_n6), .Y(
        aes_core_enc_block_n84) );
  INVX1 aes_core_enc_block_U150 ( .A(aes_core_enc_block_n239), .Y(
        aes_core_enc_block_n96) );
  INVX1 aes_core_enc_block_U149 ( .A(aes_core_enc_block_n239), .Y(
        aes_core_enc_block_n97) );
  INVX1 aes_core_enc_block_U148 ( .A(aes_core_enc_block_n239), .Y(
        aes_core_enc_block_n98) );
  INVX1 aes_core_enc_block_U147 ( .A(aes_core_enc_block_n98), .Y(
        aes_core_enc_block_n92) );
  INVX1 aes_core_enc_block_U146 ( .A(aes_core_enc_block_n709), .Y(
        aes_core_enc_block_n21) );
  CLKINVX3 aes_core_enc_block_U145 ( .A(aes_core_enc_block_n21), .Y(
        aes_core_enc_block_n20) );
  NAND2X1 aes_core_enc_block_U144 ( .A(aes_core_enc_block_n706), .B(
        aes_core_enc_block_n125), .Y(aes_core_enc_block_n233) );
  NAND2X1 aes_core_enc_block_U143 ( .A(aes_core_enc_block_n706), .B(
        aes_core_enc_block_n130), .Y(aes_core_enc_block_n468) );
  NAND2X1 aes_core_enc_block_U142 ( .A(aes_core_enc_block_n706), .B(
        aes_core_enc_block_n231), .Y(aes_core_enc_block_n948) );
  NOR3X1 aes_core_enc_block_U141 ( .A(aes_core_enc_block_n106), .B(
        aes_core_enc_block_n29), .C(aes_core_enc_block_n117), .Y(
        aes_core_enc_block_n706) );
  INVX1 aes_core_enc_block_U140 ( .A(aes_core_enc_block_n128), .Y(
        aes_core_enc_block_n127) );
  CLKINVX3 aes_core_enc_block_U139 ( .A(aes_core_enc_block_n128), .Y(
        aes_core_enc_block_n126) );
  CLKINVX3 aes_core_enc_block_U138 ( .A(aes_core_enc_block_n1), .Y(
        aes_core_enc_block_n131) );
  INVX1 aes_core_enc_block_U137 ( .A(aes_core_enc_block_n85), .Y(
        aes_core_enc_block_n75) );
  INVX1 aes_core_enc_block_U136 ( .A(aes_core_enc_block_n88), .Y(
        aes_core_enc_block_n74) );
  INVX1 aes_core_enc_block_U135 ( .A(aes_core_enc_block_n85), .Y(
        aes_core_enc_block_n81) );
  INVX1 aes_core_enc_block_U134 ( .A(aes_core_enc_block_n89), .Y(
        aes_core_enc_block_n72) );
  INVX1 aes_core_enc_block_U133 ( .A(aes_core_enc_block_n90), .Y(
        aes_core_enc_block_n70) );
  INVX1 aes_core_enc_block_U132 ( .A(aes_core_enc_block_n88), .Y(
        aes_core_enc_block_n73) );
  INVX1 aes_core_enc_block_U131 ( .A(aes_core_enc_block_n86), .Y(
        aes_core_enc_block_n79) );
  INVX1 aes_core_enc_block_U130 ( .A(aes_core_enc_block_n90), .Y(
        aes_core_enc_block_n71) );
  INVX1 aes_core_enc_block_U129 ( .A(aes_core_enc_block_n87), .Y(
        aes_core_enc_block_n76) );
  INVX1 aes_core_enc_block_U128 ( .A(aes_core_enc_block_n85), .Y(
        aes_core_enc_block_n80) );
  INVX1 aes_core_enc_block_U127 ( .A(aes_core_enc_block_n86), .Y(
        aes_core_enc_block_n78) );
  INVX1 aes_core_enc_block_U126 ( .A(aes_core_enc_block_n87), .Y(
        aes_core_enc_block_n77) );
  INVX1 aes_core_enc_block_U125 ( .A(aes_core_enc_block_n84), .Y(
        aes_core_enc_block_n82) );
  INVX1 aes_core_enc_block_U124 ( .A(aes_core_enc_block_n92), .Y(
        aes_core_enc_block_n108) );
  INVX1 aes_core_enc_block_U123 ( .A(aes_core_enc_block_n92), .Y(
        aes_core_enc_block_n107) );
  INVX1 aes_core_enc_block_U122 ( .A(aes_core_enc_block_n91), .Y(
        aes_core_enc_block_n69) );
  INVX1 aes_core_enc_block_U121 ( .A(aes_core_enc_block_n91), .Y(
        aes_core_enc_block_n68) );
  INVX1 aes_core_enc_block_U120 ( .A(aes_core_enc_block_n96), .Y(
        aes_core_enc_block_n94) );
  INVX1 aes_core_enc_block_U119 ( .A(aes_core_enc_block_n96), .Y(
        aes_core_enc_block_n95) );
  INVX1 aes_core_enc_block_U118 ( .A(aes_core_enc_block_n97), .Y(
        aes_core_enc_block_n93) );
  INVX1 aes_core_enc_block_U117 ( .A(aes_core_enc_block_n84), .Y(
        aes_core_enc_block_n83) );
  INVX1 aes_core_enc_block_U116 ( .A(aes_core_enc_block_n83), .Y(
        aes_core_enc_block_n29) );
  INVX1 aes_core_enc_block_U115 ( .A(aes_core_enc_block_n92), .Y(
        aes_core_enc_block_n106) );
  INVX1 aes_core_enc_block_U114 ( .A(aes_core_enc_block_n233), .Y(
        aes_core_enc_block_n124) );
  CLKINVX3 aes_core_enc_block_U113 ( .A(aes_core_enc_block_n124), .Y(
        aes_core_enc_block_n123) );
  INVX1 aes_core_enc_block_U112 ( .A(aes_core_enc_block_n468), .Y(
        aes_core_enc_block_n23) );
  CLKINVX3 aes_core_enc_block_U111 ( .A(aes_core_enc_block_n23), .Y(
        aes_core_enc_block_n22) );
  INVX1 aes_core_enc_block_U110 ( .A(aes_core_enc_block_n948), .Y(
        aes_core_enc_block_n19) );
  CLKINVX3 aes_core_enc_block_U109 ( .A(aes_core_enc_block_n19), .Y(
        aes_core_enc_block_n18) );
  INVX1 aes_core_enc_block_U108 ( .A(aes_core_enc_block_n230), .Y(
        aes_core_enc_block_n15) );
  INVX1 aes_core_enc_block_U107 ( .A(aes_core_enc_block_n75), .Y(
        aes_core_enc_block_n47) );
  INVX1 aes_core_enc_block_U106 ( .A(aes_core_enc_block_n81), .Y(
        aes_core_enc_block_n34) );
  INVX1 aes_core_enc_block_U105 ( .A(aes_core_enc_block_n72), .Y(
        aes_core_enc_block_n56) );
  INVX1 aes_core_enc_block_U104 ( .A(aes_core_enc_block_n70), .Y(
        aes_core_enc_block_n63) );
  INVX1 aes_core_enc_block_U103 ( .A(aes_core_enc_block_n81), .Y(
        aes_core_enc_block_n33) );
  INVX1 aes_core_enc_block_U102 ( .A(aes_core_enc_block_n73), .Y(
        aes_core_enc_block_n55) );
  INVX1 aes_core_enc_block_U101 ( .A(aes_core_enc_block_n81), .Y(
        aes_core_enc_block_n32) );
  INVX1 aes_core_enc_block_U100 ( .A(aes_core_enc_block_n73), .Y(
        aes_core_enc_block_n54) );
  INVX1 aes_core_enc_block_U99 ( .A(aes_core_enc_block_n70), .Y(
        aes_core_enc_block_n62) );
  INVX1 aes_core_enc_block_U98 ( .A(aes_core_enc_block_n79), .Y(
        aes_core_enc_block_n39) );
  INVX1 aes_core_enc_block_U97 ( .A(aes_core_enc_block_n76), .Y(
        aes_core_enc_block_n46) );
  INVX1 aes_core_enc_block_U96 ( .A(aes_core_enc_block_n74), .Y(
        aes_core_enc_block_n53) );
  INVX1 aes_core_enc_block_U95 ( .A(aes_core_enc_block_n80), .Y(
        aes_core_enc_block_n37) );
  INVX1 aes_core_enc_block_U94 ( .A(aes_core_enc_block_n76), .Y(
        aes_core_enc_block_n45) );
  INVX1 aes_core_enc_block_U93 ( .A(aes_core_enc_block_n74), .Y(
        aes_core_enc_block_n52) );
  INVX1 aes_core_enc_block_U92 ( .A(aes_core_enc_block_n80), .Y(
        aes_core_enc_block_n36) );
  INVX1 aes_core_enc_block_U91 ( .A(aes_core_enc_block_n75), .Y(
        aes_core_enc_block_n48) );
  INVX1 aes_core_enc_block_U90 ( .A(aes_core_enc_block_n75), .Y(
        aes_core_enc_block_n51) );
  INVX1 aes_core_enc_block_U89 ( .A(aes_core_enc_block_n78), .Y(
        aes_core_enc_block_n40) );
  INVX1 aes_core_enc_block_U88 ( .A(aes_core_enc_block_n77), .Y(
        aes_core_enc_block_n42) );
  INVX1 aes_core_enc_block_U87 ( .A(aes_core_enc_block_n71), .Y(
        aes_core_enc_block_n60) );
  INVX1 aes_core_enc_block_U86 ( .A(aes_core_enc_block_n76), .Y(
        aes_core_enc_block_n44) );
  INVX1 aes_core_enc_block_U85 ( .A(aes_core_enc_block_n77), .Y(
        aes_core_enc_block_n43) );
  INVX1 aes_core_enc_block_U84 ( .A(aes_core_enc_block_n71), .Y(
        aes_core_enc_block_n61) );
  INVX1 aes_core_enc_block_U83 ( .A(aes_core_enc_block_n82), .Y(
        aes_core_enc_block_n30) );
  INVX1 aes_core_enc_block_U82 ( .A(aes_core_enc_block_n79), .Y(
        aes_core_enc_block_n38) );
  INVX1 aes_core_enc_block_U81 ( .A(aes_core_enc_block_n72), .Y(
        aes_core_enc_block_n58) );
  INVX1 aes_core_enc_block_U80 ( .A(aes_core_enc_block_n72), .Y(
        aes_core_enc_block_n59) );
  INVX1 aes_core_enc_block_U79 ( .A(aes_core_enc_block_n75), .Y(
        aes_core_enc_block_n50) );
  INVX1 aes_core_enc_block_U78 ( .A(aes_core_enc_block_n75), .Y(
        aes_core_enc_block_n49) );
  INVX1 aes_core_enc_block_U77 ( .A(aes_core_enc_block_n72), .Y(
        aes_core_enc_block_n57) );
  INVX1 aes_core_enc_block_U76 ( .A(aes_core_enc_block_n80), .Y(
        aes_core_enc_block_n35) );
  INVX1 aes_core_enc_block_U75 ( .A(aes_core_enc_block_n78), .Y(
        aes_core_enc_block_n41) );
  INVX1 aes_core_enc_block_U74 ( .A(aes_core_enc_block_n82), .Y(
        aes_core_enc_block_n31) );
  INVX1 aes_core_enc_block_U73 ( .A(aes_core_enc_block_n69), .Y(
        aes_core_enc_block_n64) );
  INVX1 aes_core_enc_block_U72 ( .A(aes_core_enc_block_n68), .Y(
        aes_core_enc_block_n66) );
  INVX1 aes_core_enc_block_U71 ( .A(aes_core_enc_block_n68), .Y(
        aes_core_enc_block_n67) );
  INVX1 aes_core_enc_block_U70 ( .A(aes_core_enc_block_n69), .Y(
        aes_core_enc_block_n65) );
  INVX1 aes_core_enc_block_U69 ( .A(aes_core_enc_block_n106), .Y(
        aes_core_enc_block_n105) );
  CLKINVX3 aes_core_enc_block_U68 ( .A(aes_core_enc_block_n108), .Y(
        aes_core_enc_block_n102) );
  CLKINVX3 aes_core_enc_block_U67 ( .A(aes_core_enc_block_n107), .Y(
        aes_core_enc_block_n103) );
  CLKINVX3 aes_core_enc_block_U66 ( .A(aes_core_enc_block_n107), .Y(
        aes_core_enc_block_n104) );
  CLKINVX3 aes_core_enc_block_U65 ( .A(aes_core_enc_block_n108), .Y(
        aes_core_enc_block_n101) );
  INVX1 aes_core_enc_block_U64 ( .A(aes_core_enc_block_n95), .Y(
        aes_core_enc_block_n115) );
  INVX1 aes_core_enc_block_U63 ( .A(aes_core_enc_block_n94), .Y(
        aes_core_enc_block_n110) );
  INVX1 aes_core_enc_block_U62 ( .A(aes_core_enc_block_n95), .Y(
        aes_core_enc_block_n113) );
  INVX1 aes_core_enc_block_U61 ( .A(aes_core_enc_block_n94), .Y(
        aes_core_enc_block_n112) );
  INVX1 aes_core_enc_block_U60 ( .A(aes_core_enc_block_n94), .Y(
        aes_core_enc_block_n111) );
  INVX1 aes_core_enc_block_U59 ( .A(aes_core_enc_block_n95), .Y(
        aes_core_enc_block_n116) );
  INVX1 aes_core_enc_block_U58 ( .A(aes_core_enc_block_n95), .Y(
        aes_core_enc_block_n114) );
  INVX1 aes_core_enc_block_U57 ( .A(aes_core_enc_block_n93), .Y(
        aes_core_enc_block_n109) );
  INVX1 aes_core_enc_block_U56 ( .A(aes_core_enc_block_n2), .Y(
        aes_core_enc_block_n17) );
  INVX1 aes_core_enc_block_U55 ( .A(aes_core_enc_block_n4), .Y(
        aes_core_enc_block_n13) );
  INVX1 aes_core_enc_block_U54 ( .A(aes_core_enc_block_n4), .Y(
        aes_core_enc_block_n12) );
  INVX1 aes_core_enc_block_U53 ( .A(aes_core_enc_block_n2), .Y(
        aes_core_enc_block_n16) );
  INVX1 aes_core_enc_block_U52 ( .A(aes_core_enc_block_n3), .Y(
        aes_core_enc_block_n8) );
  INVX1 aes_core_enc_block_U51 ( .A(aes_core_enc_block_n3), .Y(
        aes_core_enc_block_n7) );
  CLKINVX3 aes_core_enc_block_U50 ( .A(aes_core_enc_block_n5), .Y(
        aes_core_enc_block_n9) );
  INVX1 aes_core_enc_block_U49 ( .A(aes_core_enc_block_n231), .Y(
        aes_core_enc_block_n11) );
  INVX1 aes_core_enc_block_U48 ( .A(aes_core_enc_block_n66), .Y(
        aes_core_enc_block_n25) );
  INVX1 aes_core_enc_block_U47 ( .A(aes_core_enc_block_n65), .Y(
        aes_core_enc_block_n24) );
  CLKINVX3 aes_core_enc_block_U46 ( .A(aes_core_enc_block_n67), .Y(
        aes_core_enc_block_n28) );
  CLKINVX3 aes_core_enc_block_U45 ( .A(aes_core_enc_block_n67), .Y(
        aes_core_enc_block_n27) );
  CLKINVX3 aes_core_enc_block_U44 ( .A(aes_core_enc_block_n66), .Y(
        aes_core_enc_block_n26) );
  INVX1 aes_core_enc_block_U43 ( .A(aes_core_enc_block_n109), .Y(
        aes_core_enc_block_n100) );
  INVX1 aes_core_enc_block_U42 ( .A(aes_core_enc_block_n109), .Y(
        aes_core_enc_block_n99) );
  OAI221X2 aes_core_enc_block_U41 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1366), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1388), .C0(aes_core_enc_block_n217), .Y(
        aes_core_enc_sboxw[20]) );
  OAI221X2 aes_core_enc_block_U40 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1437), .B0(aes_core_enc_block_n127), .B1(
        aes_core_enc_block_n1436), .C0(aes_core_enc_block_n198), .Y(
        aes_core_enc_sboxw[9]) );
  INVX8 aes_core_enc_block_U39 ( .A(aes_core_enc_round_nr[2]), .Y(
        aes_core_enc_block_n185) );
  OAI221X2 aes_core_enc_block_U38 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1376), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1385), .C0(aes_core_enc_block_n204), .Y(
        aes_core_enc_sboxw[3]) );
  INVX8 aes_core_enc_block_U37 ( .A(aes_core_enc_round_nr[1]), .Y(
        aes_core_enc_block_n184) );
  AOI22X4 aes_core_enc_block_U36 ( .A0(aes_core_enc_block_enc_ctrl_reg[0]), 
        .A1(aes_core_enc_block_n180), .B0(aes_core_enc_block_n183), .B1(
        aes_core_enc_block_n1194), .Y(aes_core_enc_block_n1193) );
  NAND2X2 aes_core_enc_block_U35 ( .A(aes_core_enc_block_n946), .B(
        aes_core_enc_block_n705), .Y(aes_core_enc_block_n230) );
  NAND2X1 aes_core_enc_block_U34 ( .A(aes_core_enc_block_n1197), .B(
        aes_core_enc_block_n1194), .Y(aes_core_enc_block_n6) );
  NOR2X4 aes_core_enc_block_U33 ( .A(aes_core_enc_block_n179), .B(
        aes_core_enc_block_n1192), .Y(aes_core_enc_block_n705) );
  NAND2X1 aes_core_enc_block_U32 ( .A(aes_core_enc_block_n705), .B(
        aes_core_enc_block_n22), .Y(aes_core_enc_block_n5) );
  NAND2X1 aes_core_enc_block_U31 ( .A(aes_core_enc_block_n705), .B(
        aes_core_enc_block_n18), .Y(aes_core_enc_block_n4) );
  NAND2X1 aes_core_enc_block_U30 ( .A(aes_core_enc_block_n705), .B(
        aes_core_enc_block_n123), .Y(aes_core_enc_block_n3) );
  NAND2X1 aes_core_enc_block_U29 ( .A(aes_core_enc_block_n705), .B(
        aes_core_enc_block_n20), .Y(aes_core_enc_block_n2) );
  OAI221X1 aes_core_enc_block_U28 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1444), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1446), .C0(aes_core_enc_block_n220), .Y(
        aes_core_enc_sboxw[18]) );
  OAI221X2 aes_core_enc_block_U27 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1347), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1398), .C0(aes_core_enc_block_n207), .Y(
        aes_core_enc_sboxw[2]) );
  INVX8 aes_core_enc_block_U26 ( .A(aes_core_enc_block_enc_ctrl_reg[0]), .Y(
        aes_core_enc_block_n181) );
  INVX8 aes_core_enc_block_U25 ( .A(aes_core_enc_block_enc_ctrl_reg[1]), .Y(
        aes_core_enc_block_n180) );
  AOI21X2 aes_core_enc_block_U24 ( .A0(aes_core_enc_block_n183), .A1(
        aes_core_enc_block_n1194), .B0(aes_core_enc_block_n1195), .Y(
        aes_core_enc_block_n1192) );
  INVX1 aes_core_enc_block_U23 ( .A(aes_core_new_sboxw[25]), .Y(
        aes_core_enc_block_n163) );
  INVX1 aes_core_enc_block_U22 ( .A(aes_core_new_sboxw[26]), .Y(
        aes_core_enc_block_n161) );
  INVX1 aes_core_enc_block_U21 ( .A(aes_core_new_sboxw[24]), .Y(
        aes_core_enc_block_n164) );
  INVX1 aes_core_enc_block_U20 ( .A(aes_core_new_sboxw[29]), .Y(
        aes_core_enc_block_n160) );
  INVX1 aes_core_enc_block_U19 ( .A(aes_core_new_sboxw[30]), .Y(
        aes_core_enc_block_n157) );
  OAI221X4 aes_core_enc_block_U18 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1374), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1364), .C0(aes_core_enc_block_n228), .Y(
        aes_core_enc_sboxw[10]) );
  INVX1 aes_core_enc_block_U17 ( .A(aes_core_enc_block_sword_ctr_reg[0]), .Y(
        aes_core_enc_block_n173) );
  INVX1 aes_core_enc_block_U16 ( .A(aes_core_enc_block_sword_ctr_reg[1]), .Y(
        aes_core_enc_block_n174) );
  OAI221X2 aes_core_enc_block_U15 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1352), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1367), .C0(aes_core_enc_block_n203), .Y(
        aes_core_enc_sboxw[4]) );
  OAI221X1 aes_core_enc_block_U14 ( .A0(aes_core_enc_block_n131), .A1(
        aes_core_enc_block_n1402), .B0(aes_core_enc_block_n126), .B1(
        aes_core_enc_block_n1387), .C0(aes_core_enc_block_n209), .Y(
        aes_core_enc_sboxw[28]) );
  OAI221X2 aes_core_enc_block_U13 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1368), .B0(aes_core_enc_block_n125), .B1(
        aes_core_enc_block_n1349), .C0(aes_core_enc_block_n226), .Y(
        aes_core_enc_sboxw[12]) );
  CLKINVX1 aes_core_enc_block_U12 ( .A(aes_core_enc_block_n197), .Y(
        aes_core_enc_block_n128) );
  AND2X1 aes_core_enc_block_U11 ( .A(aes_core_enc_block_n707), .B(
        aes_core_enc_block_n705), .Y(aes_core_enc_block_n1) );
  INVX4 aes_core_enc_block_U10 ( .A(aes_core_enc_block_n1), .Y(
        aes_core_enc_block_n130) );
  INVX12 aes_core_enc_block_U9 ( .A(aes_core_enc_block_n230), .Y(
        aes_core_enc_block_n14) );
  CLKINVX8 aes_core_enc_block_U8 ( .A(aes_core_enc_block_n231), .Y(
        aes_core_enc_block_n10) );
  NAND2X2 aes_core_enc_block_U7 ( .A(aes_core_enc_block_n1185), .B(
        aes_core_enc_block_n705), .Y(aes_core_enc_block_n231) );
  INVX1 aes_core_enc_block_U6 ( .A(aes_core_enc_round_nr[3]), .Y(
        aes_core_enc_block_n186) );
  CLKINVX3 aes_core_enc_block_U5 ( .A(aes_core_enc_block_n197), .Y(
        aes_core_enc_block_n129) );
  INVX4 aes_core_enc_block_U4 ( .A(aes_core_enc_block_n129), .Y(
        aes_core_enc_block_n125) );
  OAI221X1 aes_core_enc_block_U3 ( .A0(aes_core_enc_block_n130), .A1(
        aes_core_enc_block_n1372), .B0(aes_core_enc_block_n127), .B1(
        aes_core_enc_block_n1422), .C0(aes_core_enc_block_n199), .Y(
        aes_core_enc_sboxw[8]) );
  DFFRHQX1 aes_core_enc_block_round_ctr_reg_reg_0_ ( .D(
        aes_core_enc_block_n1342), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_round_nr[0]) );
  DFFRHQX1 aes_core_enc_block_sword_ctr_reg_reg_0_ ( .D(
        aes_core_enc_block_n1346), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_block_sword_ctr_reg[0]) );
  DFFRHQX1 aes_core_enc_block_sword_ctr_reg_reg_1_ ( .D(
        aes_core_enc_block_n1345), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_block_sword_ctr_reg[1]) );
  DFFRHQX4 aes_core_enc_block_round_ctr_reg_reg_1_ ( .D(
        aes_core_enc_block_n1341), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_round_nr[1]) );
  DFFRHQX4 aes_core_enc_block_round_ctr_reg_reg_2_ ( .D(
        aes_core_enc_block_n175), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_round_nr[2]) );
  DFFRHQX4 aes_core_enc_block_round_ctr_reg_reg_3_ ( .D(
        aes_core_enc_block_n1340), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_round_nr[3]) );
  DFFRHQX4 aes_core_enc_block_enc_ctrl_reg_reg_1_ ( .D(
        aes_core_enc_block_n1344), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_block_enc_ctrl_reg[1]) );
  DFFRHQX4 aes_core_enc_block_enc_ctrl_reg_reg_0_ ( .D(
        aes_core_enc_block_n1343), .CK(clk_48Mhz), .RN(reset_n), .Q(
        aes_core_enc_block_enc_ctrl_reg[0]) );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_27_ ( .D(
        aes_core_enc_block_n1310), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[27])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_27_ ( .D(
        aes_core_enc_block_n1278), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[59])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_27_ ( .D(
        aes_core_enc_block_n1246), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[91])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_25_ ( .D(
        aes_core_enc_block_n1248), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[89])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_24_ ( .D(
        aes_core_enc_block_n1249), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[88])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_16_ ( .D(
        aes_core_enc_block_n1321), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[16])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_19_ ( .D(
        aes_core_enc_block_n1318), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[19])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_12_ ( .D(
        aes_core_enc_block_n1325), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[12])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_16_ ( .D(
        aes_core_enc_block_n1289), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[48])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_19_ ( .D(
        aes_core_enc_block_n1286), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[51])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_11_ ( .D(
        aes_core_enc_block_n1294), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[43])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_27_ ( .D(
        aes_core_enc_block_n1215), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[123])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_11_ ( .D(
        aes_core_enc_block_n1326), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[11])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_17_ ( .D(
        aes_core_enc_block_n1256), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[81])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_16_ ( .D(
        aes_core_enc_block_n1257), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[80])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_19_ ( .D(
        aes_core_enc_block_n1254), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[83])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_20_ ( .D(
        aes_core_enc_block_n1253), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[84])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_28_ ( .D(
        aes_core_enc_block_n1245), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[92])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_17_ ( .D(
        aes_core_enc_block_n1320), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[17])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_20_ ( .D(
        aes_core_enc_block_n1317), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[20])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_4_ ( .D(
        aes_core_enc_block_n1333), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[4])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_17_ ( .D(
        aes_core_enc_block_n1288), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[49])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_20_ ( .D(
        aes_core_enc_block_n1285), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[52])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_19_ ( .D(
        aes_core_enc_block_n1223), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[115])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_16_ ( .D(
        aes_core_enc_block_n1226), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[112])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_0_ ( .D(
        aes_core_enc_block_n1338), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[96])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_25_ ( .D(
        aes_core_enc_block_n1217), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[121])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_24_ ( .D(
        aes_core_enc_block_n1218), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[120])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_28_ ( .D(
        aes_core_enc_block_n1214), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[124])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_3_ ( .D(
        aes_core_enc_block_n1334), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[3])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_0_ ( .D(
        aes_core_enc_block_n1337), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[0])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_0_ ( .D(
        aes_core_enc_block_n1305), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[32])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_3_ ( .D(
        aes_core_enc_block_n1302), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[35])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_11_ ( .D(
        aes_core_enc_block_n1231), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[107])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_9_ ( .D(
        aes_core_enc_block_n1264), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[73])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_17_ ( .D(
        aes_core_enc_block_n1225), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[113])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_13_ ( .D(
        aes_core_enc_block_n1260), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[77])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_11_ ( .D(
        aes_core_enc_block_n1262), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[75])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_20_ ( .D(
        aes_core_enc_block_n1222), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[116])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_3_ ( .D(
        aes_core_enc_block_n1239), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[99])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_3_ ( .D(
        aes_core_enc_block_n1270), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[67])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_8_ ( .D(
        aes_core_enc_block_n1265), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[72])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_12_ ( .D(
        aes_core_enc_block_n1261), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[76])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_4_ ( .D(
        aes_core_enc_block_n1269), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[68])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_1_ ( .D(
        aes_core_enc_block_n1272), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[65])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_1_ ( .D(
        aes_core_enc_block_n1336), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[1])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_1_ ( .D(
        aes_core_enc_block_n1304), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[33])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_4_ ( .D(
        aes_core_enc_block_n1301), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[36])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_9_ ( .D(
        aes_core_enc_block_n1233), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[105])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_8_ ( .D(
        aes_core_enc_block_n1234), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[104])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_12_ ( .D(
        aes_core_enc_block_n1230), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[108])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_4_ ( .D(
        aes_core_enc_block_n1238), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[100])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_1_ ( .D(
        aes_core_enc_block_n1241), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[97])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_13_ ( .D(
        aes_core_enc_block_n1229), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[109])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_26_ ( .D(
        aes_core_enc_block_n1311), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[26])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_25_ ( .D(
        aes_core_enc_block_n1312), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[25])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_24_ ( .D(
        aes_core_enc_block_n1313), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[24])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_28_ ( .D(
        aes_core_enc_block_n1309), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[28])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_26_ ( .D(
        aes_core_enc_block_n1279), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[58])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_24_ ( .D(
        aes_core_enc_block_n1281), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[56])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_29_ ( .D(
        aes_core_enc_block_n1308), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[29])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_25_ ( .D(
        aes_core_enc_block_n1280), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[57])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_29_ ( .D(
        aes_core_enc_block_n1276), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[61])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_28_ ( .D(
        aes_core_enc_block_n1277), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[60])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_26_ ( .D(
        aes_core_enc_block_n1247), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[90])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_18_ ( .D(
        aes_core_enc_block_n1319), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[18])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_18_ ( .D(
        aes_core_enc_block_n1287), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[50])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_8_ ( .D(
        aes_core_enc_block_n1297), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[40])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_10_ ( .D(
        aes_core_enc_block_n1295), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[42])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_18_ ( .D(
        aes_core_enc_block_n1255), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[82])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_21_ ( .D(
        aes_core_enc_block_n1252), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[85])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_29_ ( .D(
        aes_core_enc_block_n1244), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[93])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_21_ ( .D(
        aes_core_enc_block_n1316), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[21])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_9_ ( .D(
        aes_core_enc_block_n1328), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[9])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_13_ ( .D(
        aes_core_enc_block_n1324), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[13])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_5_ ( .D(
        aes_core_enc_block_n1332), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[5])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_21_ ( .D(
        aes_core_enc_block_n1284), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[53])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_9_ ( .D(
        aes_core_enc_block_n1296), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[41])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_18_ ( .D(
        aes_core_enc_block_n1224), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[114])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_26_ ( .D(
        aes_core_enc_block_n1216), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[122])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_10_ ( .D(
        aes_core_enc_block_n1327), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[10])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_2_ ( .D(
        aes_core_enc_block_n1335), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[2])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_2_ ( .D(
        aes_core_enc_block_n1303), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[34])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_2_ ( .D(
        aes_core_enc_block_n1240), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[98])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_21_ ( .D(
        aes_core_enc_block_n1221), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[117])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_10_ ( .D(
        aes_core_enc_block_n1263), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[74])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_5_ ( .D(
        aes_core_enc_block_n1268), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[69])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_2_ ( .D(
        aes_core_enc_block_n1271), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[66])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_29_ ( .D(
        aes_core_enc_block_n1213), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[125])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_8_ ( .D(
        aes_core_enc_block_n1329), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[8])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_12_ ( .D(
        aes_core_enc_block_n1293), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[44])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_13_ ( .D(
        aes_core_enc_block_n1292), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[45])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_5_ ( .D(
        aes_core_enc_block_n1300), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[37])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_10_ ( .D(
        aes_core_enc_block_n1232), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[106])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_5_ ( .D(
        aes_core_enc_block_n1237), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[101])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_22_ ( .D(
        aes_core_enc_block_n1251), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[86])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_30_ ( .D(
        aes_core_enc_block_n1243), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[94])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_22_ ( .D(
        aes_core_enc_block_n1315), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[22])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_6_ ( .D(
        aes_core_enc_block_n1331), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[6])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_22_ ( .D(
        aes_core_enc_block_n1283), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[54])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_22_ ( .D(
        aes_core_enc_block_n1220), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[118])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_14_ ( .D(
        aes_core_enc_block_n1259), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[78])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_6_ ( .D(
        aes_core_enc_block_n1267), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[70])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_6_ ( .D(
        aes_core_enc_block_n1236), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[102])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_14_ ( .D(
        aes_core_enc_block_n1228), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[110])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_7_ ( .D(
        aes_core_enc_block_n1330), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[7])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_7_ ( .D(
        aes_core_enc_block_n1266), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[71])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_31_ ( .D(
        aes_core_enc_block_n1242), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[95])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_7_ ( .D(
        aes_core_enc_block_n1298), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[39])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_31_ ( .D(
        aes_core_enc_block_n1306), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[31])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_30_ ( .D(
        aes_core_enc_block_n1307), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[30])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_31_ ( .D(
        aes_core_enc_block_n1274), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[63])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_30_ ( .D(
        aes_core_enc_block_n1275), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[62])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_23_ ( .D(
        aes_core_enc_block_n1250), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[87])
         );
  DFFRHQX1 aes_core_enc_block_block_w1_reg_reg_15_ ( .D(
        aes_core_enc_block_n1258), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[79])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_23_ ( .D(
        aes_core_enc_block_n1314), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[23])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_14_ ( .D(
        aes_core_enc_block_n1323), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[14])
         );
  DFFRHQX1 aes_core_enc_block_block_w3_reg_reg_15_ ( .D(
        aes_core_enc_block_n1322), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[15])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_23_ ( .D(
        aes_core_enc_block_n1282), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[55])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_7_ ( .D(
        aes_core_enc_block_n1235), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[103])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_31_ ( .D(
        aes_core_enc_block_n1211), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[127])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_30_ ( .D(
        aes_core_enc_block_n1212), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[126])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_15_ ( .D(
        aes_core_enc_block_n1290), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[47])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_14_ ( .D(
        aes_core_enc_block_n1291), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[46])
         );
  DFFRHQX1 aes_core_enc_block_block_w2_reg_reg_6_ ( .D(
        aes_core_enc_block_n1299), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[38])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_23_ ( .D(
        aes_core_enc_block_n1219), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[119])
         );
  DFFRHQX1 aes_core_enc_block_block_w0_reg_reg_15_ ( .D(
        aes_core_enc_block_n1227), .CK(clk_48Mhz), .RN(reset_n), .Q(Dout[111])
         );
  DFFSX1 aes_core_enc_block_ready_reg_reg ( .D(aes_core_enc_block_n1339), .CK(
        clk_48Mhz), .SN(reset_n), .Q(aes_core_enc_ready), .QN() );
  NAND2X1 aes_core_keymem_U2903 ( .A(aes_core_keymem_n2765), .B(
        aes_core_keymem_n24), .Y(aes_core_keymem_n838) );
  OAI2BB1X1 aes_core_keymem_U2902 ( .A0N(aes_core_keymem_key_mem_ctrl_reg[1]), 
        .A1N(aes_core_keymem_n24), .B0(aes_core_keymem_n545), .Y(
        aes_core_keymem_n543) );
  NAND3X1 aes_core_keymem_U2901 ( .A(aes_core_keymem_n17), .B(
        aes_core_keymem_n2765), .C(init), .Y(aes_core_keymem_n545) );
  NAND2X1 aes_core_keymem_U2900 ( .A(aes_core_keymem_key_mem_ctrl_reg[1]), .B(
        aes_core_keymem_n17), .Y(aes_core_keymem_n829) );
  NAND2X4 aes_core_keymem_U2899 ( .A(aes_core_keymem_key_mem_ctrl_reg[1]), .B(
        aes_core_keymem_n2763), .Y(aes_core_keymem_n22) );
  OAI2BB2X1 aes_core_keymem_U2898 ( .B0(aes_core_keymem_n2770), .B1(
        aes_core_keymem_n543), .A0N(aes_core_keymem_n543), .A1N(
        aes_core_keymem_key_mem_ctrl_reg[1]), .Y(aes_core_keymem_n841) );
  INVX1 aes_core_keymem_U2897 ( .A(aes_core_keymem_key_mem_ctrl_reg[1]), .Y(
        aes_core_keymem_n2765) );
  XNOR2X1 aes_core_keymem_U2896 ( .A(aes_core_keymem_rcon_reg[0]), .B(
        aes_core_keymem_rcon_reg[7]), .Y(aes_core_keymem_n833) );
  NOR2X1 aes_core_keymem_U2895 ( .A(aes_core_keymem_n833), .B(
        aes_core_keymem_n829), .Y(aes_core_keymem_n2384) );
  XNOR2X1 aes_core_keymem_U2894 ( .A(aes_core_keymem_rcon_reg[3]), .B(
        aes_core_keymem_rcon_reg[7]), .Y(aes_core_keymem_n831) );
  NOR2X1 aes_core_keymem_U2893 ( .A(aes_core_keymem_n831), .B(
        aes_core_keymem_n829), .Y(aes_core_keymem_n2381) );
  OAI22X1 aes_core_keymem_U2892 ( .A0(aes_core_keymem_n2767), .A1(
        aes_core_keymem_n834), .B0(aes_core_keymem_round_ctr_reg[0]), .B1(
        aes_core_keymem_n829), .Y(aes_core_keymem_n2386) );
  INVX1 aes_core_keymem_U2891 ( .A(aes_core_key_ready), .Y(
        aes_core_keymem_n2770) );
  INVX1 aes_core_keymem_U2890 ( .A(init), .Y(aes_core_keymem_n2773) );
  AND2X2 aes_core_keymem_U2889 ( .A(aes_core_keymem_rcon_reg[4]), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2380) );
  AND2X2 aes_core_keymem_U2888 ( .A(aes_core_keymem_rcon_reg[5]), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2379) );
  XNOR2X1 aes_core_keymem_U2887 ( .A(aes_core_keymem_rcon_reg[2]), .B(
        aes_core_keymem_rcon_reg[7]), .Y(aes_core_keymem_n832) );
  NAND2X1 aes_core_keymem_U2886 ( .A(aes_core_keymem_n832), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2382) );
  NAND2BX1 aes_core_keymem_U2885 ( .AN(aes_core_keymem_rcon_reg[6]), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2378) );
  NAND2BX1 aes_core_keymem_U2884 ( .AN(aes_core_keymem_rcon_reg[1]), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2383) );
  NAND2BX1 aes_core_keymem_U2883 ( .AN(aes_core_keymem_rcon_reg[7]), .B(
        aes_core_keymem_n2762), .Y(aes_core_keymem_n2385) );
  OAI21X1 aes_core_keymem_U2882 ( .A0(aes_core_keymem_round_ctr_reg[0]), .A1(
        aes_core_keymem_n829), .B0(aes_core_keymem_n834), .Y(
        aes_core_keymem_n836) );
  AND2X1 aes_core_keymem_U2881 ( .A(aes_core_enc_round_nr[3]), .B(
        aes_core_enc_round_nr[1]), .Y(aes_core_keymem_n23) );
  AND3X1 aes_core_keymem_U2880 ( .A(aes_core_enc_round_nr[0]), .B(
        aes_core_enc_round_nr[1]), .C(aes_core_enc_round_nr[2]), .Y(
        aes_core_keymem_n26) );
  INVX1 aes_core_keymem_U2879 ( .A(aes_core_keymem_n825), .Y(
        aes_core_keymem_n2766) );
  OAI32X1 aes_core_keymem_U2878 ( .A0(aes_core_keymem_n2766), .A1(
        aes_core_keymem_round_ctr_reg[2]), .A2(aes_core_keymem_n829), .B0(
        aes_core_keymem_n837), .B1(aes_core_keymem_n2769), .Y(
        aes_core_keymem_n2387) );
  NOR2X1 aes_core_keymem_U2877 ( .A(aes_core_keymem_round_ctr_reg[2]), .B(
        aes_core_keymem_round_ctr_reg[3]), .Y(aes_core_keymem_n828) );
  AOI22X1 aes_core_keymem_U2876 ( .A0(aes_core_keymem_n836), .A1(
        aes_core_keymem_round_ctr_reg[1]), .B0(aes_core_keymem_n2762), .B1(
        aes_core_keymem_n824), .Y(aes_core_keymem_n835) );
  INVX1 aes_core_keymem_U2875 ( .A(aes_core_keymem_n835), .Y(
        aes_core_keymem_n2761) );
  AOI222X1 aes_core_keymem_U2874 ( .A0(aes_core_keymem_key_mem[351]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[95]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[223]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n51) );
  AOI222X1 aes_core_keymem_U2873 ( .A0(aes_core_keymem_key_mem[863]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[607]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[735]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n52) );
  AOI22X1 aes_core_keymem_U2872 ( .A0(aes_core_keymem_key_mem[1247]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1375]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n49) );
  NAND4X1 aes_core_keymem_U2871 ( .A(aes_core_keymem_n49), .B(
        aes_core_keymem_n50), .C(aes_core_keymem_n51), .D(aes_core_keymem_n52), 
        .Y(aes_core_round_key[95]) );
  AOI222X1 aes_core_keymem_U2870 ( .A0(aes_core_keymem_key_mem[349]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[93]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[221]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n59) );
  AOI222X1 aes_core_keymem_U2869 ( .A0(aes_core_keymem_key_mem[861]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[605]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[733]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n60) );
  AOI22X1 aes_core_keymem_U2868 ( .A0(aes_core_keymem_key_mem[1245]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1373]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n57) );
  NAND4X1 aes_core_keymem_U2867 ( .A(aes_core_keymem_n57), .B(
        aes_core_keymem_n58), .C(aes_core_keymem_n59), .D(aes_core_keymem_n60), 
        .Y(aes_core_round_key[93]) );
  AOI222X1 aes_core_keymem_U2866 ( .A0(aes_core_keymem_key_mem[350]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[94]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[222]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n55) );
  AOI222X1 aes_core_keymem_U2865 ( .A0(aes_core_keymem_key_mem[862]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[606]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[734]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n56) );
  AOI22X1 aes_core_keymem_U2864 ( .A0(aes_core_keymem_key_mem[1246]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1374]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n53) );
  NAND4X1 aes_core_keymem_U2863 ( .A(aes_core_keymem_n53), .B(
        aes_core_keymem_n54), .C(aes_core_keymem_n55), .D(aes_core_keymem_n56), 
        .Y(aes_core_round_key[94]) );
  AOI222X1 aes_core_keymem_U2862 ( .A0(aes_core_keymem_key_mem[380]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[124]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[252]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n431) );
  AOI222X1 aes_core_keymem_U2861 ( .A0(aes_core_keymem_key_mem[892]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[636]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[764]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n432) );
  AOI22X1 aes_core_keymem_U2860 ( .A0(aes_core_keymem_key_mem[1276]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1404]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n429) );
  NAND4X1 aes_core_keymem_U2859 ( .A(aes_core_keymem_n429), .B(
        aes_core_keymem_n430), .C(aes_core_keymem_n431), .D(
        aes_core_keymem_n432), .Y(aes_core_round_key[124]) );
  AOI222X1 aes_core_keymem_U2858 ( .A0(aes_core_keymem_key_mem[284]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[28]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[156]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n347) );
  AOI222X1 aes_core_keymem_U2857 ( .A0(aes_core_keymem_key_mem[796]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[540]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[668]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n348) );
  AOI22X1 aes_core_keymem_U2856 ( .A0(aes_core_keymem_key_mem[1180]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1308]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n345) );
  NAND4X1 aes_core_keymem_U2855 ( .A(aes_core_keymem_n345), .B(
        aes_core_keymem_n346), .C(aes_core_keymem_n347), .D(
        aes_core_keymem_n348), .Y(aes_core_round_key[28]) );
  AOI222X1 aes_core_keymem_U2854 ( .A0(aes_core_keymem_key_mem[316]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[60]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[188]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n203) );
  AOI222X1 aes_core_keymem_U2853 ( .A0(aes_core_keymem_key_mem[828]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[572]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[700]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n204) );
  AOI22X1 aes_core_keymem_U2852 ( .A0(aes_core_keymem_key_mem[1212]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1340]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n201) );
  NAND4X1 aes_core_keymem_U2851 ( .A(aes_core_keymem_n201), .B(
        aes_core_keymem_n202), .C(aes_core_keymem_n203), .D(
        aes_core_keymem_n204), .Y(aes_core_round_key[60]) );
  AOI222X1 aes_core_keymem_U2850 ( .A0(aes_core_keymem_key_mem[348]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[92]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[220]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n63) );
  AOI222X1 aes_core_keymem_U2849 ( .A0(aes_core_keymem_key_mem[860]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[604]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[732]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n64) );
  AOI22X1 aes_core_keymem_U2848 ( .A0(aes_core_keymem_key_mem[1244]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1372]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n61) );
  NAND4X1 aes_core_keymem_U2847 ( .A(aes_core_keymem_n61), .B(
        aes_core_keymem_n62), .C(aes_core_keymem_n63), .D(aes_core_keymem_n64), 
        .Y(aes_core_round_key[92]) );
  AOI222X1 aes_core_keymem_U2846 ( .A0(aes_core_keymem_key_mem[345]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[89]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[217]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n79) );
  AOI222X1 aes_core_keymem_U2845 ( .A0(aes_core_keymem_key_mem[857]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[601]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[729]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n80) );
  AOI22X1 aes_core_keymem_U2844 ( .A0(aes_core_keymem_key_mem[1241]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1369]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n77) );
  NAND4X1 aes_core_keymem_U2843 ( .A(aes_core_keymem_n77), .B(
        aes_core_keymem_n78), .C(aes_core_keymem_n79), .D(aes_core_keymem_n80), 
        .Y(aes_core_round_key[89]) );
  AOI222X1 aes_core_keymem_U2842 ( .A0(aes_core_keymem_key_mem[377]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[121]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[249]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n443) );
  AOI222X1 aes_core_keymem_U2841 ( .A0(aes_core_keymem_key_mem[889]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[633]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[761]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n444) );
  AOI22X1 aes_core_keymem_U2840 ( .A0(aes_core_keymem_key_mem[1273]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1401]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n441) );
  NAND4X1 aes_core_keymem_U2839 ( .A(aes_core_keymem_n441), .B(
        aes_core_keymem_n442), .C(aes_core_keymem_n443), .D(
        aes_core_keymem_n444), .Y(aes_core_round_key[121]) );
  AOI222X1 aes_core_keymem_U2838 ( .A0(aes_core_keymem_key_mem[281]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[25]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[153]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n359) );
  AOI222X1 aes_core_keymem_U2837 ( .A0(aes_core_keymem_key_mem[793]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[537]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[665]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n360) );
  AOI22X1 aes_core_keymem_U2836 ( .A0(aes_core_keymem_key_mem[1177]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1305]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n357) );
  NAND4X1 aes_core_keymem_U2835 ( .A(aes_core_keymem_n357), .B(
        aes_core_keymem_n358), .C(aes_core_keymem_n359), .D(
        aes_core_keymem_n360), .Y(aes_core_round_key[25]) );
  AOI222X1 aes_core_keymem_U2834 ( .A0(aes_core_keymem_key_mem[313]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[57]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[185]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n219) );
  AOI222X1 aes_core_keymem_U2833 ( .A0(aes_core_keymem_key_mem[825]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[569]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[697]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n220) );
  AOI22X1 aes_core_keymem_U2832 ( .A0(aes_core_keymem_key_mem[1209]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1337]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n217) );
  NAND4X1 aes_core_keymem_U2831 ( .A(aes_core_keymem_n217), .B(
        aes_core_keymem_n218), .C(aes_core_keymem_n219), .D(
        aes_core_keymem_n220), .Y(aes_core_round_key[57]) );
  AOI222X1 aes_core_keymem_U2830 ( .A0(aes_core_keymem_key_mem[379]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[123]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[251]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n435) );
  AOI222X1 aes_core_keymem_U2829 ( .A0(aes_core_keymem_key_mem[891]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[635]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[763]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n436) );
  AOI22X1 aes_core_keymem_U2828 ( .A0(aes_core_keymem_key_mem[1275]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1403]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n433) );
  NAND4X1 aes_core_keymem_U2827 ( .A(aes_core_keymem_n433), .B(
        aes_core_keymem_n434), .C(aes_core_keymem_n435), .D(
        aes_core_keymem_n436), .Y(aes_core_round_key[123]) );
  AOI222X1 aes_core_keymem_U2826 ( .A0(aes_core_keymem_key_mem[283]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[27]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[155]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n351) );
  AOI222X1 aes_core_keymem_U2825 ( .A0(aes_core_keymem_key_mem[795]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[539]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[667]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n352) );
  AOI22X1 aes_core_keymem_U2824 ( .A0(aes_core_keymem_key_mem[1179]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1307]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n349) );
  NAND4X1 aes_core_keymem_U2823 ( .A(aes_core_keymem_n349), .B(
        aes_core_keymem_n350), .C(aes_core_keymem_n351), .D(
        aes_core_keymem_n352), .Y(aes_core_round_key[27]) );
  AOI222X1 aes_core_keymem_U2822 ( .A0(aes_core_keymem_key_mem[347]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[91]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[219]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n67) );
  AOI222X1 aes_core_keymem_U2821 ( .A0(aes_core_keymem_key_mem[859]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[603]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[731]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n68) );
  AOI22X1 aes_core_keymem_U2820 ( .A0(aes_core_keymem_key_mem[1243]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1371]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n65) );
  NAND4X1 aes_core_keymem_U2819 ( .A(aes_core_keymem_n65), .B(
        aes_core_keymem_n66), .C(aes_core_keymem_n67), .D(aes_core_keymem_n68), 
        .Y(aes_core_round_key[91]) );
  AOI222X1 aes_core_keymem_U2818 ( .A0(aes_core_keymem_key_mem[315]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[59]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[187]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n211) );
  AOI222X1 aes_core_keymem_U2817 ( .A0(aes_core_keymem_key_mem[827]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[571]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[699]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n212) );
  AOI22X1 aes_core_keymem_U2816 ( .A0(aes_core_keymem_key_mem[1211]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1339]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n209) );
  NAND4X1 aes_core_keymem_U2815 ( .A(aes_core_keymem_n209), .B(
        aes_core_keymem_n210), .C(aes_core_keymem_n211), .D(
        aes_core_keymem_n212), .Y(aes_core_round_key[59]) );
  AOI222X1 aes_core_keymem_U2814 ( .A0(aes_core_keymem_key_mem[285]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[29]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[157]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n343) );
  AOI222X1 aes_core_keymem_U2813 ( .A0(aes_core_keymem_key_mem[797]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[541]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[669]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n344) );
  AOI22X1 aes_core_keymem_U2812 ( .A0(aes_core_keymem_key_mem[1181]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1309]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n341) );
  NAND4X1 aes_core_keymem_U2811 ( .A(aes_core_keymem_n341), .B(
        aes_core_keymem_n342), .C(aes_core_keymem_n343), .D(
        aes_core_keymem_n344), .Y(aes_core_round_key[29]) );
  AOI222X1 aes_core_keymem_U2810 ( .A0(aes_core_keymem_key_mem[286]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[30]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[158]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n335) );
  AOI222X1 aes_core_keymem_U2809 ( .A0(aes_core_keymem_key_mem[798]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[542]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[670]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n336) );
  AOI22X1 aes_core_keymem_U2808 ( .A0(aes_core_keymem_key_mem[1182]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1310]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n333) );
  NAND4X1 aes_core_keymem_U2807 ( .A(aes_core_keymem_n333), .B(
        aes_core_keymem_n334), .C(aes_core_keymem_n335), .D(
        aes_core_keymem_n336), .Y(aes_core_round_key[30]) );
  AOI222X1 aes_core_keymem_U2806 ( .A0(aes_core_keymem_key_mem[287]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[31]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[159]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n331) );
  AOI222X1 aes_core_keymem_U2805 ( .A0(aes_core_keymem_key_mem[799]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[543]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[671]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n332) );
  AOI22X1 aes_core_keymem_U2804 ( .A0(aes_core_keymem_key_mem[1183]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1311]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n329) );
  NAND4X1 aes_core_keymem_U2803 ( .A(aes_core_keymem_n329), .B(
        aes_core_keymem_n330), .C(aes_core_keymem_n331), .D(
        aes_core_keymem_n332), .Y(aes_core_round_key[31]) );
  AOI222X1 aes_core_keymem_U2802 ( .A0(aes_core_keymem_key_mem[317]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[61]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[189]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n199) );
  AOI222X1 aes_core_keymem_U2801 ( .A0(aes_core_keymem_key_mem[829]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[573]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[701]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n200) );
  AOI22X1 aes_core_keymem_U2800 ( .A0(aes_core_keymem_key_mem[1213]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1341]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n197) );
  NAND4X1 aes_core_keymem_U2799 ( .A(aes_core_keymem_n197), .B(
        aes_core_keymem_n198), .C(aes_core_keymem_n199), .D(
        aes_core_keymem_n200), .Y(aes_core_round_key[61]) );
  AOI222X1 aes_core_keymem_U2798 ( .A0(aes_core_keymem_key_mem[318]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[62]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[190]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n195) );
  AOI222X1 aes_core_keymem_U2797 ( .A0(aes_core_keymem_key_mem[830]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[574]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[702]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n196) );
  AOI22X1 aes_core_keymem_U2796 ( .A0(aes_core_keymem_key_mem[1214]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1342]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n193) );
  NAND4X1 aes_core_keymem_U2795 ( .A(aes_core_keymem_n193), .B(
        aes_core_keymem_n194), .C(aes_core_keymem_n195), .D(
        aes_core_keymem_n196), .Y(aes_core_round_key[62]) );
  AOI222X1 aes_core_keymem_U2794 ( .A0(aes_core_keymem_key_mem[319]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[63]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[191]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n191) );
  AOI222X1 aes_core_keymem_U2793 ( .A0(aes_core_keymem_key_mem[831]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[575]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[703]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n192) );
  AOI22X1 aes_core_keymem_U2792 ( .A0(aes_core_keymem_key_mem[1215]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1343]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n189) );
  NAND4X1 aes_core_keymem_U2791 ( .A(aes_core_keymem_n189), .B(
        aes_core_keymem_n190), .C(aes_core_keymem_n191), .D(
        aes_core_keymem_n192), .Y(aes_core_round_key[63]) );
  AOI222X1 aes_core_keymem_U2790 ( .A0(aes_core_keymem_key_mem[312]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[56]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[184]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n223) );
  AOI222X1 aes_core_keymem_U2789 ( .A0(aes_core_keymem_key_mem[824]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[568]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[696]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n224) );
  AOI22X1 aes_core_keymem_U2788 ( .A0(aes_core_keymem_key_mem[1208]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1336]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n221) );
  NAND4X1 aes_core_keymem_U2787 ( .A(aes_core_keymem_n221), .B(
        aes_core_keymem_n222), .C(aes_core_keymem_n223), .D(
        aes_core_keymem_n224), .Y(aes_core_round_key[56]) );
  AOI222X1 aes_core_keymem_U2786 ( .A0(aes_core_keymem_key_mem[381]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[125]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[253]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n427) );
  AOI222X1 aes_core_keymem_U2785 ( .A0(aes_core_keymem_key_mem[893]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[637]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[765]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n428) );
  AOI22X1 aes_core_keymem_U2784 ( .A0(aes_core_keymem_key_mem[1277]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1405]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n425) );
  NAND4X1 aes_core_keymem_U2783 ( .A(aes_core_keymem_n425), .B(
        aes_core_keymem_n426), .C(aes_core_keymem_n427), .D(
        aes_core_keymem_n428), .Y(aes_core_round_key[125]) );
  AOI222X1 aes_core_keymem_U2782 ( .A0(aes_core_keymem_key_mem[382]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[126]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[254]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n423) );
  AOI222X1 aes_core_keymem_U2781 ( .A0(aes_core_keymem_key_mem[894]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[638]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[766]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n424) );
  AOI22X1 aes_core_keymem_U2780 ( .A0(aes_core_keymem_key_mem[1278]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1406]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n421) );
  NAND4X1 aes_core_keymem_U2779 ( .A(aes_core_keymem_n421), .B(
        aes_core_keymem_n422), .C(aes_core_keymem_n423), .D(
        aes_core_keymem_n424), .Y(aes_core_round_key[126]) );
  AOI222X1 aes_core_keymem_U2778 ( .A0(aes_core_keymem_key_mem[383]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[127]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[255]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n419) );
  AOI222X1 aes_core_keymem_U2777 ( .A0(aes_core_keymem_key_mem[895]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[639]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[767]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n420) );
  AOI22X1 aes_core_keymem_U2776 ( .A0(aes_core_keymem_key_mem[1279]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1407]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n417) );
  NAND4X1 aes_core_keymem_U2775 ( .A(aes_core_keymem_n417), .B(
        aes_core_keymem_n418), .C(aes_core_keymem_n419), .D(
        aes_core_keymem_n420), .Y(aes_core_round_key[127]) );
  AOI222X1 aes_core_keymem_U2774 ( .A0(aes_core_keymem_key_mem[376]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[120]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[248]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n447) );
  AOI222X1 aes_core_keymem_U2773 ( .A0(aes_core_keymem_key_mem[888]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[632]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[760]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n448) );
  AOI22X1 aes_core_keymem_U2772 ( .A0(aes_core_keymem_key_mem[1272]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1400]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n445) );
  NAND4X1 aes_core_keymem_U2771 ( .A(aes_core_keymem_n445), .B(
        aes_core_keymem_n446), .C(aes_core_keymem_n447), .D(
        aes_core_keymem_n448), .Y(aes_core_round_key[120]) );
  AOI222X1 aes_core_keymem_U2770 ( .A0(aes_core_keymem_key_mem[280]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[24]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[152]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n363) );
  AOI222X1 aes_core_keymem_U2769 ( .A0(aes_core_keymem_key_mem[792]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[536]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[664]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n364) );
  AOI22X1 aes_core_keymem_U2768 ( .A0(aes_core_keymem_key_mem[1176]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1304]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n361) );
  NAND4X1 aes_core_keymem_U2767 ( .A(aes_core_keymem_n361), .B(
        aes_core_keymem_n362), .C(aes_core_keymem_n363), .D(
        aes_core_keymem_n364), .Y(aes_core_round_key[24]) );
  AOI222X1 aes_core_keymem_U2766 ( .A0(aes_core_keymem_key_mem[344]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[88]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[216]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n83) );
  AOI222X1 aes_core_keymem_U2765 ( .A0(aes_core_keymem_key_mem[856]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[600]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[728]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n84) );
  AOI22X1 aes_core_keymem_U2764 ( .A0(aes_core_keymem_key_mem[1240]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1368]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n81) );
  NAND4X1 aes_core_keymem_U2763 ( .A(aes_core_keymem_n81), .B(
        aes_core_keymem_n82), .C(aes_core_keymem_n83), .D(aes_core_keymem_n84), 
        .Y(aes_core_round_key[88]) );
  AOI222X1 aes_core_keymem_U2762 ( .A0(aes_core_keymem_key_mem[314]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[58]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[186]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n215) );
  AOI222X1 aes_core_keymem_U2761 ( .A0(aes_core_keymem_key_mem[826]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[570]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[698]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n216) );
  AOI22X1 aes_core_keymem_U2760 ( .A0(aes_core_keymem_key_mem[1210]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1338]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n213) );
  NAND4X1 aes_core_keymem_U2759 ( .A(aes_core_keymem_n213), .B(
        aes_core_keymem_n214), .C(aes_core_keymem_n215), .D(
        aes_core_keymem_n216), .Y(aes_core_round_key[58]) );
  AOI222X1 aes_core_keymem_U2758 ( .A0(aes_core_keymem_key_mem[346]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[90]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[218]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n71) );
  AOI222X1 aes_core_keymem_U2757 ( .A0(aes_core_keymem_key_mem[858]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[602]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[730]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n72) );
  AOI22X1 aes_core_keymem_U2756 ( .A0(aes_core_keymem_key_mem[1242]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1370]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n69) );
  NAND4X1 aes_core_keymem_U2755 ( .A(aes_core_keymem_n69), .B(
        aes_core_keymem_n70), .C(aes_core_keymem_n71), .D(aes_core_keymem_n72), 
        .Y(aes_core_round_key[90]) );
  AOI222X1 aes_core_keymem_U2754 ( .A0(aes_core_keymem_key_mem[378]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[122]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[250]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n439) );
  AOI222X1 aes_core_keymem_U2753 ( .A0(aes_core_keymem_key_mem[890]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[634]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[762]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n440) );
  AOI22X1 aes_core_keymem_U2752 ( .A0(aes_core_keymem_key_mem[1274]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1402]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n437) );
  NAND4X1 aes_core_keymem_U2751 ( .A(aes_core_keymem_n437), .B(
        aes_core_keymem_n438), .C(aes_core_keymem_n439), .D(
        aes_core_keymem_n440), .Y(aes_core_round_key[122]) );
  AOI222X1 aes_core_keymem_U2750 ( .A0(aes_core_keymem_key_mem[282]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[26]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[154]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n355) );
  AOI222X1 aes_core_keymem_U2749 ( .A0(aes_core_keymem_key_mem[794]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[538]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[666]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n356) );
  AOI22X1 aes_core_keymem_U2748 ( .A0(aes_core_keymem_key_mem[1178]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1306]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n353) );
  NAND4X1 aes_core_keymem_U2747 ( .A(aes_core_keymem_n353), .B(
        aes_core_keymem_n354), .C(aes_core_keymem_n355), .D(
        aes_core_keymem_n356), .Y(aes_core_round_key[26]) );
  NOR2X1 aes_core_keymem_U2746 ( .A(aes_core_enc_round_nr[2]), .B(
        aes_core_enc_round_nr[3]), .Y(aes_core_keymem_n542) );
  NOR2X1 aes_core_keymem_U2745 ( .A(aes_core_enc_round_nr[0]), .B(
        aes_core_enc_round_nr[1]), .Y(aes_core_keymem_n541) );
  INVX1 aes_core_keymem_U2744 ( .A(aes_core_enc_round_nr[0]), .Y(
        aes_core_keymem_n2771) );
  AOI222X1 aes_core_keymem_U2743 ( .A0(aes_core_keymem_key_mem[352]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[96]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[224]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n47) );
  AOI222X1 aes_core_keymem_U2742 ( .A0(aes_core_keymem_key_mem[864]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[608]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[736]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n48) );
  AOI22X1 aes_core_keymem_U2741 ( .A0(aes_core_keymem_key_mem[1248]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1376]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n45) );
  NAND4X1 aes_core_keymem_U2740 ( .A(aes_core_keymem_n45), .B(
        aes_core_keymem_n46), .C(aes_core_keymem_n47), .D(aes_core_keymem_n48), 
        .Y(aes_core_round_key[96]) );
  AOI222X1 aes_core_keymem_U2739 ( .A0(aes_core_keymem_key_mem[353]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[97]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[225]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n43) );
  AOI222X1 aes_core_keymem_U2738 ( .A0(aes_core_keymem_key_mem[865]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[609]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[737]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n44) );
  AOI22X1 aes_core_keymem_U2737 ( .A0(aes_core_keymem_key_mem[1249]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1377]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n41) );
  NAND4X1 aes_core_keymem_U2736 ( .A(aes_core_keymem_n41), .B(
        aes_core_keymem_n42), .C(aes_core_keymem_n43), .D(aes_core_keymem_n44), 
        .Y(aes_core_round_key[97]) );
  AOI222X1 aes_core_keymem_U2735 ( .A0(aes_core_keymem_key_mem[265]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[9]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[137]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n20) );
  AOI222X1 aes_core_keymem_U2734 ( .A0(aes_core_keymem_key_mem[777]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[521]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[649]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n21) );
  AOI22X1 aes_core_keymem_U2733 ( .A0(aes_core_keymem_key_mem[1161]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1289]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n18) );
  NAND4X1 aes_core_keymem_U2732 ( .A(aes_core_keymem_n18), .B(
        aes_core_keymem_n19), .C(aes_core_keymem_n20), .D(aes_core_keymem_n21), 
        .Y(aes_core_round_key[9]) );
  AOI222X1 aes_core_keymem_U2731 ( .A0(aes_core_keymem_key_mem[355]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[99]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[227]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n35) );
  AOI222X1 aes_core_keymem_U2730 ( .A0(aes_core_keymem_key_mem[867]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[611]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[739]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n36) );
  AOI22X1 aes_core_keymem_U2729 ( .A0(aes_core_keymem_key_mem[1251]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1379]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n33) );
  NAND4X1 aes_core_keymem_U2728 ( .A(aes_core_keymem_n33), .B(
        aes_core_keymem_n34), .C(aes_core_keymem_n35), .D(aes_core_keymem_n36), 
        .Y(aes_core_round_key[99]) );
  AOI222X1 aes_core_keymem_U2727 ( .A0(aes_core_keymem_key_mem[354]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[98]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[226]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n39) );
  AOI222X1 aes_core_keymem_U2726 ( .A0(aes_core_keymem_key_mem[866]), .A1(
        aes_core_keymem_n2760), .B0(aes_core_keymem_key_mem[610]), .B1(
        aes_core_keymem_n23), .C0(aes_core_keymem_key_mem[738]), .C1(
        aes_core_keymem_n2738), .Y(aes_core_keymem_n40) );
  AOI22X1 aes_core_keymem_U2725 ( .A0(aes_core_keymem_key_mem[1250]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1378]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n37) );
  NAND4X1 aes_core_keymem_U2724 ( .A(aes_core_keymem_n37), .B(
        aes_core_keymem_n38), .C(aes_core_keymem_n39), .D(aes_core_keymem_n40), 
        .Y(aes_core_round_key[98]) );
  AOI222X1 aes_core_keymem_U2723 ( .A0(aes_core_keymem_key_mem[321]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[65]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[193]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n183) );
  AOI222X1 aes_core_keymem_U2722 ( .A0(aes_core_keymem_key_mem[833]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[577]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[705]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n184) );
  AOI22X1 aes_core_keymem_U2721 ( .A0(aes_core_keymem_key_mem[1217]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1345]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n181) );
  NAND4X1 aes_core_keymem_U2720 ( .A(aes_core_keymem_n181), .B(
        aes_core_keymem_n182), .C(aes_core_keymem_n183), .D(
        aes_core_keymem_n184), .Y(aes_core_round_key[65]) );
  AOI222X1 aes_core_keymem_U2719 ( .A0(aes_core_keymem_key_mem[298]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[42]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[170]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n283) );
  AOI222X1 aes_core_keymem_U2718 ( .A0(aes_core_keymem_key_mem[810]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[554]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[682]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n284) );
  AOI22X1 aes_core_keymem_U2717 ( .A0(aes_core_keymem_key_mem[1194]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1322]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n281) );
  NAND4X1 aes_core_keymem_U2716 ( .A(aes_core_keymem_n281), .B(
        aes_core_keymem_n282), .C(aes_core_keymem_n283), .D(
        aes_core_keymem_n284), .Y(aes_core_round_key[42]) );
  AOI222X1 aes_core_keymem_U2715 ( .A0(aes_core_keymem_key_mem[363]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[107]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[235]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n507) );
  AOI222X1 aes_core_keymem_U2714 ( .A0(aes_core_keymem_key_mem[875]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[619]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[747]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n508) );
  AOI22X1 aes_core_keymem_U2713 ( .A0(aes_core_keymem_key_mem[1259]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1387]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n505) );
  NAND4X1 aes_core_keymem_U2712 ( .A(aes_core_keymem_n505), .B(
        aes_core_keymem_n506), .C(aes_core_keymem_n507), .D(
        aes_core_keymem_n508), .Y(aes_core_round_key[107]) );
  AOI222X1 aes_core_keymem_U2711 ( .A0(aes_core_keymem_key_mem[291]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[35]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[163]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n315) );
  AOI222X1 aes_core_keymem_U2710 ( .A0(aes_core_keymem_key_mem[803]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[547]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[675]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n316) );
  AOI22X1 aes_core_keymem_U2709 ( .A0(aes_core_keymem_key_mem[1187]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1315]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n313) );
  NAND4X1 aes_core_keymem_U2708 ( .A(aes_core_keymem_n313), .B(
        aes_core_keymem_n314), .C(aes_core_keymem_n315), .D(
        aes_core_keymem_n316), .Y(aes_core_round_key[35]) );
  AOI222X1 aes_core_keymem_U2707 ( .A0(aes_core_keymem_key_mem[260]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[4]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[132]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n251) );
  AOI222X1 aes_core_keymem_U2706 ( .A0(aes_core_keymem_key_mem[772]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[516]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[644]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n252) );
  AOI22X1 aes_core_keymem_U2705 ( .A0(aes_core_keymem_key_mem[1156]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1284]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n249) );
  NAND4X1 aes_core_keymem_U2704 ( .A(aes_core_keymem_n249), .B(
        aes_core_keymem_n250), .C(aes_core_keymem_n251), .D(
        aes_core_keymem_n252), .Y(aes_core_round_key[4]) );
  AOI222X1 aes_core_keymem_U2703 ( .A0(aes_core_keymem_key_mem[365]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[109]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[237]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n499) );
  AOI222X1 aes_core_keymem_U2702 ( .A0(aes_core_keymem_key_mem[877]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[621]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[749]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n500) );
  AOI22X1 aes_core_keymem_U2701 ( .A0(aes_core_keymem_key_mem[1261]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1389]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n497) );
  NAND4X1 aes_core_keymem_U2700 ( .A(aes_core_keymem_n497), .B(
        aes_core_keymem_n498), .C(aes_core_keymem_n499), .D(
        aes_core_keymem_n500), .Y(aes_core_round_key[109]) );
  AOI222X1 aes_core_keymem_U2699 ( .A0(aes_core_keymem_key_mem[293]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[37]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[165]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n307) );
  AOI222X1 aes_core_keymem_U2698 ( .A0(aes_core_keymem_key_mem[805]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[549]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[677]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n308) );
  AOI22X1 aes_core_keymem_U2697 ( .A0(aes_core_keymem_key_mem[1189]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1317]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n305) );
  NAND4X1 aes_core_keymem_U2696 ( .A(aes_core_keymem_n305), .B(
        aes_core_keymem_n306), .C(aes_core_keymem_n307), .D(
        aes_core_keymem_n308), .Y(aes_core_round_key[37]) );
  AOI222X1 aes_core_keymem_U2695 ( .A0(aes_core_keymem_key_mem[261]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[5]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[133]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n207) );
  AOI222X1 aes_core_keymem_U2694 ( .A0(aes_core_keymem_key_mem[773]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[517]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[645]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n208) );
  AOI22X1 aes_core_keymem_U2693 ( .A0(aes_core_keymem_key_mem[1157]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1285]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n205) );
  NAND4X1 aes_core_keymem_U2692 ( .A(aes_core_keymem_n205), .B(
        aes_core_keymem_n206), .C(aes_core_keymem_n207), .D(
        aes_core_keymem_n208), .Y(aes_core_round_key[5]) );
  AOI222X1 aes_core_keymem_U2691 ( .A0(aes_core_keymem_key_mem[366]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[110]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[238]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n491) );
  AOI222X1 aes_core_keymem_U2690 ( .A0(aes_core_keymem_key_mem[878]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[622]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[750]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n492) );
  AOI22X1 aes_core_keymem_U2689 ( .A0(aes_core_keymem_key_mem[1262]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1390]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n489) );
  NAND4X1 aes_core_keymem_U2688 ( .A(aes_core_keymem_n489), .B(
        aes_core_keymem_n490), .C(aes_core_keymem_n491), .D(
        aes_core_keymem_n492), .Y(aes_core_round_key[110]) );
  AOI222X1 aes_core_keymem_U2687 ( .A0(aes_core_keymem_key_mem[294]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[38]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[166]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n303) );
  AOI222X1 aes_core_keymem_U2686 ( .A0(aes_core_keymem_key_mem[806]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[550]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[678]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n304) );
  AOI22X1 aes_core_keymem_U2685 ( .A0(aes_core_keymem_key_mem[1190]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1318]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n301) );
  NAND4X1 aes_core_keymem_U2684 ( .A(aes_core_keymem_n301), .B(
        aes_core_keymem_n302), .C(aes_core_keymem_n303), .D(
        aes_core_keymem_n304), .Y(aes_core_round_key[38]) );
  AOI222X1 aes_core_keymem_U2683 ( .A0(aes_core_keymem_key_mem[262]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[6]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[134]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n163) );
  AOI222X1 aes_core_keymem_U2682 ( .A0(aes_core_keymem_key_mem[774]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[518]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[646]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n164) );
  AOI22X1 aes_core_keymem_U2681 ( .A0(aes_core_keymem_key_mem[1158]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1286]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n161) );
  NAND4X1 aes_core_keymem_U2680 ( .A(aes_core_keymem_n161), .B(
        aes_core_keymem_n162), .C(aes_core_keymem_n163), .D(
        aes_core_keymem_n164), .Y(aes_core_round_key[6]) );
  AOI222X1 aes_core_keymem_U2679 ( .A0(aes_core_keymem_key_mem[367]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[111]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[239]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n487) );
  AOI222X1 aes_core_keymem_U2678 ( .A0(aes_core_keymem_key_mem[879]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[623]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[751]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n488) );
  AOI22X1 aes_core_keymem_U2677 ( .A0(aes_core_keymem_key_mem[1263]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1391]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n485) );
  NAND4X1 aes_core_keymem_U2676 ( .A(aes_core_keymem_n485), .B(
        aes_core_keymem_n486), .C(aes_core_keymem_n487), .D(
        aes_core_keymem_n488), .Y(aes_core_round_key[111]) );
  AOI222X1 aes_core_keymem_U2675 ( .A0(aes_core_keymem_key_mem[295]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[39]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[167]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n299) );
  AOI222X1 aes_core_keymem_U2674 ( .A0(aes_core_keymem_key_mem[807]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[551]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[679]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n300) );
  AOI22X1 aes_core_keymem_U2673 ( .A0(aes_core_keymem_key_mem[1191]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1319]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n297) );
  NAND4X1 aes_core_keymem_U2672 ( .A(aes_core_keymem_n297), .B(
        aes_core_keymem_n298), .C(aes_core_keymem_n299), .D(
        aes_core_keymem_n300), .Y(aes_core_round_key[39]) );
  AOI222X1 aes_core_keymem_U2671 ( .A0(aes_core_keymem_key_mem[256]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[0]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[128]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n539) );
  AOI222X1 aes_core_keymem_U2670 ( .A0(aes_core_keymem_key_mem[768]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[512]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[640]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n540) );
  AOI22X1 aes_core_keymem_U2669 ( .A0(aes_core_keymem_key_mem[1152]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1280]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n537) );
  NAND4X1 aes_core_keymem_U2668 ( .A(aes_core_keymem_n537), .B(
        aes_core_keymem_n538), .C(aes_core_keymem_n539), .D(
        aes_core_keymem_n540), .Y(aes_core_round_key[0]) );
  AOI222X1 aes_core_keymem_U2667 ( .A0(aes_core_keymem_key_mem[322]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[66]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[194]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n179) );
  AOI222X1 aes_core_keymem_U2666 ( .A0(aes_core_keymem_key_mem[834]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[578]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[706]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n180) );
  AOI22X1 aes_core_keymem_U2665 ( .A0(aes_core_keymem_key_mem[1218]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1346]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n177) );
  NAND4X1 aes_core_keymem_U2664 ( .A(aes_core_keymem_n177), .B(
        aes_core_keymem_n178), .C(aes_core_keymem_n179), .D(
        aes_core_keymem_n180), .Y(aes_core_round_key[66]) );
  AOI222X1 aes_core_keymem_U2663 ( .A0(aes_core_keymem_key_mem[299]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[43]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[171]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n279) );
  AOI222X1 aes_core_keymem_U2662 ( .A0(aes_core_keymem_key_mem[811]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[555]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[683]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n280) );
  AOI22X1 aes_core_keymem_U2661 ( .A0(aes_core_keymem_key_mem[1195]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1323]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n277) );
  NAND4X1 aes_core_keymem_U2660 ( .A(aes_core_keymem_n277), .B(
        aes_core_keymem_n278), .C(aes_core_keymem_n279), .D(
        aes_core_keymem_n280), .Y(aes_core_round_key[43]) );
  AOI222X1 aes_core_keymem_U2659 ( .A0(aes_core_keymem_key_mem[364]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[108]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[236]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n503) );
  AOI222X1 aes_core_keymem_U2658 ( .A0(aes_core_keymem_key_mem[876]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[620]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[748]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n504) );
  AOI22X1 aes_core_keymem_U2657 ( .A0(aes_core_keymem_key_mem[1260]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1388]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n501) );
  NAND4X1 aes_core_keymem_U2656 ( .A(aes_core_keymem_n501), .B(
        aes_core_keymem_n502), .C(aes_core_keymem_n503), .D(
        aes_core_keymem_n504), .Y(aes_core_round_key[108]) );
  AOI222X1 aes_core_keymem_U2655 ( .A0(aes_core_keymem_key_mem[292]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[36]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[164]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n311) );
  AOI222X1 aes_core_keymem_U2654 ( .A0(aes_core_keymem_key_mem[804]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[548]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[676]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n312) );
  AOI22X1 aes_core_keymem_U2653 ( .A0(aes_core_keymem_key_mem[1188]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1316]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n309) );
  NAND4X1 aes_core_keymem_U2652 ( .A(aes_core_keymem_n309), .B(
        aes_core_keymem_n310), .C(aes_core_keymem_n311), .D(
        aes_core_keymem_n312), .Y(aes_core_round_key[36]) );
  AOI222X1 aes_core_keymem_U2651 ( .A0(aes_core_keymem_key_mem[268]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[12]), .B1(
        aes_core_keymem_n2715), .C0(aes_core_keymem_key_mem[140]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n415) );
  AOI222X1 aes_core_keymem_U2650 ( .A0(aes_core_keymem_key_mem[780]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[524]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[652]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n416) );
  AOI22X1 aes_core_keymem_U2649 ( .A0(aes_core_keymem_key_mem[1164]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1292]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n413) );
  NAND4X1 aes_core_keymem_U2648 ( .A(aes_core_keymem_n413), .B(
        aes_core_keymem_n414), .C(aes_core_keymem_n415), .D(
        aes_core_keymem_n416), .Y(aes_core_round_key[12]) );
  AOI222X1 aes_core_keymem_U2647 ( .A0(aes_core_keymem_key_mem[324]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[68]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[196]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n171) );
  AOI222X1 aes_core_keymem_U2646 ( .A0(aes_core_keymem_key_mem[836]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[580]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[708]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n172) );
  AOI22X1 aes_core_keymem_U2645 ( .A0(aes_core_keymem_key_mem[1220]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1348]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n169) );
  NAND4X1 aes_core_keymem_U2644 ( .A(aes_core_keymem_n169), .B(
        aes_core_keymem_n170), .C(aes_core_keymem_n171), .D(
        aes_core_keymem_n172), .Y(aes_core_round_key[68]) );
  AOI222X1 aes_core_keymem_U2643 ( .A0(aes_core_keymem_key_mem[301]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[45]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[173]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n271) );
  AOI222X1 aes_core_keymem_U2642 ( .A0(aes_core_keymem_key_mem[813]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[557]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[685]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n272) );
  AOI22X1 aes_core_keymem_U2641 ( .A0(aes_core_keymem_key_mem[1197]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1325]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n269) );
  NAND4X1 aes_core_keymem_U2640 ( .A(aes_core_keymem_n269), .B(
        aes_core_keymem_n270), .C(aes_core_keymem_n271), .D(
        aes_core_keymem_n272), .Y(aes_core_round_key[45]) );
  AOI222X1 aes_core_keymem_U2639 ( .A0(aes_core_keymem_key_mem[357]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[101]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[229]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n531) );
  AOI222X1 aes_core_keymem_U2638 ( .A0(aes_core_keymem_key_mem[869]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[613]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[741]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n532) );
  AOI22X1 aes_core_keymem_U2637 ( .A0(aes_core_keymem_key_mem[1253]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1381]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n529) );
  NAND4X1 aes_core_keymem_U2636 ( .A(aes_core_keymem_n529), .B(
        aes_core_keymem_n530), .C(aes_core_keymem_n531), .D(
        aes_core_keymem_n532), .Y(aes_core_round_key[101]) );
  AOI222X1 aes_core_keymem_U2635 ( .A0(aes_core_keymem_key_mem[325]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[69]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[197]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n167) );
  AOI222X1 aes_core_keymem_U2634 ( .A0(aes_core_keymem_key_mem[837]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[581]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[709]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n168) );
  AOI22X1 aes_core_keymem_U2633 ( .A0(aes_core_keymem_key_mem[1221]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1349]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n165) );
  NAND4X1 aes_core_keymem_U2632 ( .A(aes_core_keymem_n165), .B(
        aes_core_keymem_n166), .C(aes_core_keymem_n167), .D(
        aes_core_keymem_n168), .Y(aes_core_round_key[69]) );
  AOI222X1 aes_core_keymem_U2631 ( .A0(aes_core_keymem_key_mem[302]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[46]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[174]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n267) );
  AOI222X1 aes_core_keymem_U2630 ( .A0(aes_core_keymem_key_mem[814]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[558]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[686]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n268) );
  AOI22X1 aes_core_keymem_U2629 ( .A0(aes_core_keymem_key_mem[1198]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1326]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n265) );
  NAND4X1 aes_core_keymem_U2628 ( .A(aes_core_keymem_n265), .B(
        aes_core_keymem_n266), .C(aes_core_keymem_n267), .D(
        aes_core_keymem_n268), .Y(aes_core_round_key[46]) );
  AOI222X1 aes_core_keymem_U2627 ( .A0(aes_core_keymem_key_mem[358]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[102]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[230]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n527) );
  AOI222X1 aes_core_keymem_U2626 ( .A0(aes_core_keymem_key_mem[870]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[614]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[742]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n528) );
  AOI22X1 aes_core_keymem_U2625 ( .A0(aes_core_keymem_key_mem[1254]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1382]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n525) );
  NAND4X1 aes_core_keymem_U2624 ( .A(aes_core_keymem_n525), .B(
        aes_core_keymem_n526), .C(aes_core_keymem_n527), .D(
        aes_core_keymem_n528), .Y(aes_core_round_key[102]) );
  AOI222X1 aes_core_keymem_U2623 ( .A0(aes_core_keymem_key_mem[326]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[70]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[198]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n159) );
  AOI222X1 aes_core_keymem_U2622 ( .A0(aes_core_keymem_key_mem[838]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[582]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[710]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n160) );
  AOI22X1 aes_core_keymem_U2621 ( .A0(aes_core_keymem_key_mem[1222]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1350]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n157) );
  NAND4X1 aes_core_keymem_U2620 ( .A(aes_core_keymem_n157), .B(
        aes_core_keymem_n158), .C(aes_core_keymem_n159), .D(
        aes_core_keymem_n160), .Y(aes_core_round_key[70]) );
  AOI222X1 aes_core_keymem_U2619 ( .A0(aes_core_keymem_key_mem[303]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[47]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[175]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n263) );
  AOI222X1 aes_core_keymem_U2618 ( .A0(aes_core_keymem_key_mem[815]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[559]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[687]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n264) );
  AOI22X1 aes_core_keymem_U2617 ( .A0(aes_core_keymem_key_mem[1199]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1327]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n261) );
  NAND4X1 aes_core_keymem_U2616 ( .A(aes_core_keymem_n261), .B(
        aes_core_keymem_n262), .C(aes_core_keymem_n263), .D(
        aes_core_keymem_n264), .Y(aes_core_round_key[47]) );
  AOI222X1 aes_core_keymem_U2615 ( .A0(aes_core_keymem_key_mem[359]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[103]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[231]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n523) );
  AOI222X1 aes_core_keymem_U2614 ( .A0(aes_core_keymem_key_mem[871]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[615]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[743]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n524) );
  AOI22X1 aes_core_keymem_U2613 ( .A0(aes_core_keymem_key_mem[1255]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1383]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n521) );
  NAND4X1 aes_core_keymem_U2612 ( .A(aes_core_keymem_n521), .B(
        aes_core_keymem_n522), .C(aes_core_keymem_n523), .D(
        aes_core_keymem_n524), .Y(aes_core_round_key[103]) );
  AOI222X1 aes_core_keymem_U2611 ( .A0(aes_core_keymem_key_mem[320]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[64]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[192]), .C1(
        aes_core_keymem_n27), .Y(aes_core_keymem_n187) );
  AOI222X1 aes_core_keymem_U2610 ( .A0(aes_core_keymem_key_mem[832]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[576]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[704]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n188) );
  AOI22X1 aes_core_keymem_U2609 ( .A0(aes_core_keymem_key_mem[1216]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1344]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n185) );
  NAND4X1 aes_core_keymem_U2608 ( .A(aes_core_keymem_n185), .B(
        aes_core_keymem_n186), .C(aes_core_keymem_n187), .D(
        aes_core_keymem_n188), .Y(aes_core_round_key[64]) );
  AOI222X1 aes_core_keymem_U2607 ( .A0(aes_core_keymem_key_mem[297]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[41]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[169]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n287) );
  AOI222X1 aes_core_keymem_U2606 ( .A0(aes_core_keymem_key_mem[809]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[553]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[681]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n288) );
  AOI22X1 aes_core_keymem_U2605 ( .A0(aes_core_keymem_key_mem[1193]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1321]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n285) );
  NAND4X1 aes_core_keymem_U2604 ( .A(aes_core_keymem_n285), .B(
        aes_core_keymem_n286), .C(aes_core_keymem_n287), .D(
        aes_core_keymem_n288), .Y(aes_core_round_key[41]) );
  AOI222X1 aes_core_keymem_U2603 ( .A0(aes_core_keymem_key_mem[362]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[106]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[234]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n511) );
  AOI222X1 aes_core_keymem_U2602 ( .A0(aes_core_keymem_key_mem[874]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[618]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[746]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n512) );
  AOI22X1 aes_core_keymem_U2601 ( .A0(aes_core_keymem_key_mem[1258]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1386]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n509) );
  NAND4X1 aes_core_keymem_U2600 ( .A(aes_core_keymem_n509), .B(
        aes_core_keymem_n510), .C(aes_core_keymem_n511), .D(
        aes_core_keymem_n512), .Y(aes_core_round_key[106]) );
  AOI222X1 aes_core_keymem_U2599 ( .A0(aes_core_keymem_key_mem[307]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[51]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[179]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n243) );
  AOI222X1 aes_core_keymem_U2598 ( .A0(aes_core_keymem_key_mem[819]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[563]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[691]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n244) );
  AOI22X1 aes_core_keymem_U2597 ( .A0(aes_core_keymem_key_mem[1203]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1331]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n241) );
  NAND4X1 aes_core_keymem_U2596 ( .A(aes_core_keymem_n241), .B(
        aes_core_keymem_n242), .C(aes_core_keymem_n243), .D(
        aes_core_keymem_n244), .Y(aes_core_round_key[51]) );
  AOI222X1 aes_core_keymem_U2595 ( .A0(aes_core_keymem_key_mem[340]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[84]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[212]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n99) );
  AOI222X1 aes_core_keymem_U2594 ( .A0(aes_core_keymem_key_mem[852]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[596]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[724]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n100) );
  AOI22X1 aes_core_keymem_U2593 ( .A0(aes_core_keymem_key_mem[1236]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1364]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n97) );
  NAND4X1 aes_core_keymem_U2592 ( .A(aes_core_keymem_n97), .B(
        aes_core_keymem_n98), .C(aes_core_keymem_n99), .D(aes_core_keymem_n100), .Y(aes_core_round_key[84]) );
  AOI222X1 aes_core_keymem_U2591 ( .A0(aes_core_keymem_key_mem[356]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[100]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[228]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n535) );
  AOI222X1 aes_core_keymem_U2590 ( .A0(aes_core_keymem_key_mem[868]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[612]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[740]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n536) );
  AOI22X1 aes_core_keymem_U2589 ( .A0(aes_core_keymem_key_mem[1252]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1380]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n533) );
  NAND4X1 aes_core_keymem_U2588 ( .A(aes_core_keymem_n533), .B(
        aes_core_keymem_n534), .C(aes_core_keymem_n535), .D(
        aes_core_keymem_n536), .Y(aes_core_round_key[100]) );
  AOI222X1 aes_core_keymem_U2587 ( .A0(aes_core_keymem_key_mem[332]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[76]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[204]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n135) );
  AOI222X1 aes_core_keymem_U2586 ( .A0(aes_core_keymem_key_mem[844]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[588]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[716]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n136) );
  AOI22X1 aes_core_keymem_U2585 ( .A0(aes_core_keymem_key_mem[1228]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1356]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n133) );
  NAND4X1 aes_core_keymem_U2584 ( .A(aes_core_keymem_n133), .B(
        aes_core_keymem_n134), .C(aes_core_keymem_n135), .D(
        aes_core_keymem_n136), .Y(aes_core_round_key[76]) );
  AOI222X1 aes_core_keymem_U2583 ( .A0(aes_core_keymem_key_mem[269]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[13]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[141]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n411) );
  AOI222X1 aes_core_keymem_U2582 ( .A0(aes_core_keymem_key_mem[781]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[525]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[653]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n412) );
  AOI22X1 aes_core_keymem_U2581 ( .A0(aes_core_keymem_key_mem[1165]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1293]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n409) );
  NAND4X1 aes_core_keymem_U2580 ( .A(aes_core_keymem_n409), .B(
        aes_core_keymem_n410), .C(aes_core_keymem_n411), .D(
        aes_core_keymem_n412), .Y(aes_core_round_key[13]) );
  AOI222X1 aes_core_keymem_U2579 ( .A0(aes_core_keymem_key_mem[334]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[78]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[206]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n127) );
  AOI222X1 aes_core_keymem_U2578 ( .A0(aes_core_keymem_key_mem[846]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[590]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[718]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n128) );
  AOI22X1 aes_core_keymem_U2577 ( .A0(aes_core_keymem_key_mem[1230]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1358]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n125) );
  NAND4X1 aes_core_keymem_U2576 ( .A(aes_core_keymem_n125), .B(
        aes_core_keymem_n126), .C(aes_core_keymem_n127), .D(
        aes_core_keymem_n128), .Y(aes_core_round_key[78]) );
  AOI222X1 aes_core_keymem_U2575 ( .A0(aes_core_keymem_key_mem[271]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[15]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[143]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n403) );
  AOI222X1 aes_core_keymem_U2574 ( .A0(aes_core_keymem_key_mem[783]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[527]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[655]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n404) );
  AOI22X1 aes_core_keymem_U2573 ( .A0(aes_core_keymem_key_mem[1167]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1295]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n401) );
  NAND4X1 aes_core_keymem_U2572 ( .A(aes_core_keymem_n401), .B(
        aes_core_keymem_n402), .C(aes_core_keymem_n403), .D(
        aes_core_keymem_n404), .Y(aes_core_round_key[15]) );
  AOI222X1 aes_core_keymem_U2571 ( .A0(aes_core_keymem_key_mem[328]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[72]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[200]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n151) );
  AOI222X1 aes_core_keymem_U2570 ( .A0(aes_core_keymem_key_mem[840]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[584]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[712]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n152) );
  AOI22X1 aes_core_keymem_U2569 ( .A0(aes_core_keymem_key_mem[1224]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1352]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n149) );
  NAND4X1 aes_core_keymem_U2568 ( .A(aes_core_keymem_n149), .B(
        aes_core_keymem_n150), .C(aes_core_keymem_n151), .D(
        aes_core_keymem_n152), .Y(aes_core_round_key[72]) );
  AOI222X1 aes_core_keymem_U2567 ( .A0(aes_core_keymem_key_mem[330]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[74]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[202]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n143) );
  AOI222X1 aes_core_keymem_U2566 ( .A0(aes_core_keymem_key_mem[842]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[586]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[714]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n144) );
  AOI22X1 aes_core_keymem_U2565 ( .A0(aes_core_keymem_key_mem[1226]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1354]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n141) );
  NAND4X1 aes_core_keymem_U2564 ( .A(aes_core_keymem_n141), .B(
        aes_core_keymem_n142), .C(aes_core_keymem_n143), .D(
        aes_core_keymem_n144), .Y(aes_core_round_key[74]) );
  AOI222X1 aes_core_keymem_U2563 ( .A0(aes_core_keymem_key_mem[267]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[11]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[139]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n451) );
  AOI222X1 aes_core_keymem_U2562 ( .A0(aes_core_keymem_key_mem[779]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[523]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[651]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n452) );
  AOI22X1 aes_core_keymem_U2561 ( .A0(aes_core_keymem_key_mem[1163]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1291]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n449) );
  NAND4X1 aes_core_keymem_U2560 ( .A(aes_core_keymem_n449), .B(
        aes_core_keymem_n450), .C(aes_core_keymem_n451), .D(
        aes_core_keymem_n452), .Y(aes_core_round_key[11]) );
  AOI222X1 aes_core_keymem_U2559 ( .A0(aes_core_keymem_key_mem[323]), .A1(
        aes_core_keymem_n2723), .B0(aes_core_keymem_key_mem[67]), .B1(
        aes_core_keymem_n2712), .C0(aes_core_keymem_key_mem[195]), .C1(
        aes_core_keymem_n2704), .Y(aes_core_keymem_n175) );
  AOI222X1 aes_core_keymem_U2558 ( .A0(aes_core_keymem_key_mem[835]), .A1(
        aes_core_keymem_n2757), .B0(aes_core_keymem_key_mem[579]), .B1(
        aes_core_keymem_n2746), .C0(aes_core_keymem_key_mem[707]), .C1(
        aes_core_keymem_n2735), .Y(aes_core_keymem_n176) );
  AOI22X1 aes_core_keymem_U2557 ( .A0(aes_core_keymem_key_mem[1219]), .A1(
        aes_core_keymem_n2658), .B0(aes_core_keymem_key_mem[1347]), .B1(
        aes_core_keymem_n2648), .Y(aes_core_keymem_n173) );
  NAND4X1 aes_core_keymem_U2556 ( .A(aes_core_keymem_n173), .B(
        aes_core_keymem_n174), .C(aes_core_keymem_n175), .D(
        aes_core_keymem_n176), .Y(aes_core_round_key[67]) );
  AOI222X1 aes_core_keymem_U2555 ( .A0(aes_core_keymem_key_mem[300]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[44]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[172]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n275) );
  AOI222X1 aes_core_keymem_U2554 ( .A0(aes_core_keymem_key_mem[812]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[556]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[684]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n276) );
  AOI22X1 aes_core_keymem_U2553 ( .A0(aes_core_keymem_key_mem[1196]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1324]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n273) );
  NAND4X1 aes_core_keymem_U2552 ( .A(aes_core_keymem_n273), .B(
        aes_core_keymem_n274), .C(aes_core_keymem_n275), .D(
        aes_core_keymem_n276), .Y(aes_core_round_key[44]) );
  AOI222X1 aes_core_keymem_U2551 ( .A0(aes_core_keymem_key_mem[373]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[117]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[245]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n463) );
  AOI222X1 aes_core_keymem_U2550 ( .A0(aes_core_keymem_key_mem[885]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[629]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[757]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n464) );
  AOI22X1 aes_core_keymem_U2549 ( .A0(aes_core_keymem_key_mem[1269]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1397]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n461) );
  NAND4X1 aes_core_keymem_U2548 ( .A(aes_core_keymem_n461), .B(
        aes_core_keymem_n462), .C(aes_core_keymem_n463), .D(
        aes_core_keymem_n464), .Y(aes_core_round_key[117]) );
  AOI222X1 aes_core_keymem_U2547 ( .A0(aes_core_keymem_key_mem[270]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[14]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[142]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n407) );
  AOI222X1 aes_core_keymem_U2546 ( .A0(aes_core_keymem_key_mem[782]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[526]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[654]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n408) );
  AOI22X1 aes_core_keymem_U2545 ( .A0(aes_core_keymem_key_mem[1166]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1294]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n405) );
  NAND4X1 aes_core_keymem_U2544 ( .A(aes_core_keymem_n405), .B(
        aes_core_keymem_n406), .C(aes_core_keymem_n407), .D(
        aes_core_keymem_n408), .Y(aes_core_round_key[14]) );
  AOI222X1 aes_core_keymem_U2543 ( .A0(aes_core_keymem_key_mem[335]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[79]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[207]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n123) );
  AOI222X1 aes_core_keymem_U2542 ( .A0(aes_core_keymem_key_mem[847]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[591]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[719]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n124) );
  AOI22X1 aes_core_keymem_U2541 ( .A0(aes_core_keymem_key_mem[1231]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1359]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n121) );
  NAND4X1 aes_core_keymem_U2540 ( .A(aes_core_keymem_n121), .B(
        aes_core_keymem_n122), .C(aes_core_keymem_n123), .D(
        aes_core_keymem_n124), .Y(aes_core_round_key[79]) );
  AOI222X1 aes_core_keymem_U2539 ( .A0(aes_core_keymem_key_mem[263]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[7]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[135]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n119) );
  AOI222X1 aes_core_keymem_U2538 ( .A0(aes_core_keymem_key_mem[775]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[519]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[647]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n120) );
  AOI22X1 aes_core_keymem_U2537 ( .A0(aes_core_keymem_key_mem[1159]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1287]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n117) );
  NAND4X1 aes_core_keymem_U2536 ( .A(aes_core_keymem_n117), .B(
        aes_core_keymem_n118), .C(aes_core_keymem_n119), .D(
        aes_core_keymem_n120), .Y(aes_core_round_key[7]) );
  AOI222X1 aes_core_keymem_U2535 ( .A0(aes_core_keymem_key_mem[339]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[83]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[211]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n103) );
  AOI222X1 aes_core_keymem_U2534 ( .A0(aes_core_keymem_key_mem[851]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[595]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[723]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n104) );
  AOI22X1 aes_core_keymem_U2533 ( .A0(aes_core_keymem_key_mem[1235]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1363]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n101) );
  NAND4X1 aes_core_keymem_U2532 ( .A(aes_core_keymem_n101), .B(
        aes_core_keymem_n102), .C(aes_core_keymem_n103), .D(
        aes_core_keymem_n104), .Y(aes_core_round_key[83]) );
  AOI222X1 aes_core_keymem_U2531 ( .A0(aes_core_keymem_key_mem[372]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[116]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[244]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n467) );
  AOI222X1 aes_core_keymem_U2530 ( .A0(aes_core_keymem_key_mem[884]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[628]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[756]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n468) );
  AOI22X1 aes_core_keymem_U2529 ( .A0(aes_core_keymem_key_mem[1268]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1396]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n465) );
  NAND4X1 aes_core_keymem_U2528 ( .A(aes_core_keymem_n465), .B(
        aes_core_keymem_n466), .C(aes_core_keymem_n467), .D(
        aes_core_keymem_n468), .Y(aes_core_round_key[116]) );
  AOI222X1 aes_core_keymem_U2527 ( .A0(aes_core_keymem_key_mem[276]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[20]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[148]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n379) );
  AOI222X1 aes_core_keymem_U2526 ( .A0(aes_core_keymem_key_mem[788]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[532]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[660]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n380) );
  AOI22X1 aes_core_keymem_U2525 ( .A0(aes_core_keymem_key_mem[1172]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1300]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n377) );
  NAND4X1 aes_core_keymem_U2524 ( .A(aes_core_keymem_n377), .B(
        aes_core_keymem_n378), .C(aes_core_keymem_n379), .D(
        aes_core_keymem_n380), .Y(aes_core_round_key[20]) );
  AOI222X1 aes_core_keymem_U2523 ( .A0(aes_core_keymem_key_mem[288]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[32]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[160]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n327) );
  AOI222X1 aes_core_keymem_U2522 ( .A0(aes_core_keymem_key_mem[800]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[544]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[672]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n328) );
  AOI22X1 aes_core_keymem_U2521 ( .A0(aes_core_keymem_key_mem[1184]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1312]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n325) );
  NAND4X1 aes_core_keymem_U2520 ( .A(aes_core_keymem_n325), .B(
        aes_core_keymem_n326), .C(aes_core_keymem_n327), .D(
        aes_core_keymem_n328), .Y(aes_core_round_key[32]) );
  AOI222X1 aes_core_keymem_U2518 ( .A0(aes_core_keymem_key_mem[257]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[1]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[129]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n383) );
  AOI222X1 aes_core_keymem_U2517 ( .A0(aes_core_keymem_key_mem[769]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[513]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[641]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n384) );
  AOI22X1 aes_core_keymem_U2516 ( .A0(aes_core_keymem_key_mem[1153]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1281]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n381) );
  NAND4X1 aes_core_keymem_U2514 ( .A(aes_core_keymem_n381), .B(
        aes_core_keymem_n382), .C(aes_core_keymem_n383), .D(
        aes_core_keymem_n384), .Y(aes_core_round_key[1]) );
  AOI222X1 aes_core_keymem_U2513 ( .A0(aes_core_keymem_key_mem[331]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[75]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[203]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n139) );
  AOI222X1 aes_core_keymem_U2512 ( .A0(aes_core_keymem_key_mem[843]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[587]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[715]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n140) );
  AOI22X1 aes_core_keymem_U2511 ( .A0(aes_core_keymem_key_mem[1227]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1355]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n137) );
  NAND4X1 aes_core_keymem_U2510 ( .A(aes_core_keymem_n137), .B(
        aes_core_keymem_n138), .C(aes_core_keymem_n139), .D(
        aes_core_keymem_n140), .Y(aes_core_round_key[75]) );
  AOI222X1 aes_core_keymem_U2509 ( .A0(aes_core_keymem_key_mem[275]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[19]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[147]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n387) );
  AOI222X1 aes_core_keymem_U2508 ( .A0(aes_core_keymem_key_mem[787]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[531]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[659]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n388) );
  AOI22X1 aes_core_keymem_U2507 ( .A0(aes_core_keymem_key_mem[1171]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1299]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n385) );
  NAND4X1 aes_core_keymem_U2506 ( .A(aes_core_keymem_n385), .B(
        aes_core_keymem_n386), .C(aes_core_keymem_n387), .D(
        aes_core_keymem_n388), .Y(aes_core_round_key[19]) );
  AOI222X1 aes_core_keymem_U2505 ( .A0(aes_core_keymem_key_mem[308]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[52]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[180]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n239) );
  AOI222X1 aes_core_keymem_U2504 ( .A0(aes_core_keymem_key_mem[820]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[564]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[692]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n240) );
  AOI22X1 aes_core_keymem_U2503 ( .A0(aes_core_keymem_key_mem[1204]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1332]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n237) );
  NAND4X1 aes_core_keymem_U2502 ( .A(aes_core_keymem_n237), .B(
        aes_core_keymem_n238), .C(aes_core_keymem_n239), .D(
        aes_core_keymem_n240), .Y(aes_core_round_key[52]) );
  AOI222X1 aes_core_keymem_U2501 ( .A0(aes_core_keymem_key_mem[333]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[77]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[205]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n131) );
  AOI222X1 aes_core_keymem_U2500 ( .A0(aes_core_keymem_key_mem[845]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[589]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[717]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n132) );
  AOI22X1 aes_core_keymem_U2499 ( .A0(aes_core_keymem_key_mem[1229]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1357]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n129) );
  NAND4X1 aes_core_keymem_U2498 ( .A(aes_core_keymem_n129), .B(
        aes_core_keymem_n130), .C(aes_core_keymem_n131), .D(
        aes_core_keymem_n132), .Y(aes_core_round_key[77]) );
  AOI222X1 aes_core_keymem_U2497 ( .A0(aes_core_keymem_key_mem[277]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[21]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[149]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n375) );
  AOI222X1 aes_core_keymem_U2496 ( .A0(aes_core_keymem_key_mem[789]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[533]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[661]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n376) );
  AOI22X1 aes_core_keymem_U2495 ( .A0(aes_core_keymem_key_mem[1173]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1301]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n373) );
  NAND4X1 aes_core_keymem_U2494 ( .A(aes_core_keymem_n373), .B(
        aes_core_keymem_n374), .C(aes_core_keymem_n375), .D(
        aes_core_keymem_n376), .Y(aes_core_round_key[21]) );
  AOI222X1 aes_core_keymem_U2493 ( .A0(aes_core_keymem_key_mem[309]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[53]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[181]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n235) );
  AOI222X1 aes_core_keymem_U2492 ( .A0(aes_core_keymem_key_mem[821]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[565]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[693]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n236) );
  AOI22X1 aes_core_keymem_U2491 ( .A0(aes_core_keymem_key_mem[1205]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1333]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n233) );
  NAND4X1 aes_core_keymem_U2490 ( .A(aes_core_keymem_n233), .B(
        aes_core_keymem_n234), .C(aes_core_keymem_n235), .D(
        aes_core_keymem_n236), .Y(aes_core_round_key[53]) );
  AOI222X1 aes_core_keymem_U2489 ( .A0(aes_core_keymem_key_mem[341]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[85]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[213]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n95) );
  AOI222X1 aes_core_keymem_U2488 ( .A0(aes_core_keymem_key_mem[853]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[597]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[725]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n96) );
  AOI22X1 aes_core_keymem_U2487 ( .A0(aes_core_keymem_key_mem[1237]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1365]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n93) );
  NAND4X1 aes_core_keymem_U2486 ( .A(aes_core_keymem_n93), .B(
        aes_core_keymem_n94), .C(aes_core_keymem_n95), .D(aes_core_keymem_n96), 
        .Y(aes_core_round_key[85]) );
  AOI222X1 aes_core_keymem_U2485 ( .A0(aes_core_keymem_key_mem[374]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[118]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[246]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n459) );
  AOI222X1 aes_core_keymem_U2484 ( .A0(aes_core_keymem_key_mem[886]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[630]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[758]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n460) );
  AOI22X1 aes_core_keymem_U2483 ( .A0(aes_core_keymem_key_mem[1270]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1398]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n457) );
  NAND4X1 aes_core_keymem_U2482 ( .A(aes_core_keymem_n457), .B(
        aes_core_keymem_n458), .C(aes_core_keymem_n459), .D(
        aes_core_keymem_n460), .Y(aes_core_round_key[118]) );
  AOI222X1 aes_core_keymem_U2481 ( .A0(aes_core_keymem_key_mem[278]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[22]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[150]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n371) );
  AOI222X1 aes_core_keymem_U2480 ( .A0(aes_core_keymem_key_mem[790]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[534]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[662]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n372) );
  AOI22X1 aes_core_keymem_U2479 ( .A0(aes_core_keymem_key_mem[1174]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1302]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n369) );
  NAND4X1 aes_core_keymem_U2478 ( .A(aes_core_keymem_n369), .B(
        aes_core_keymem_n370), .C(aes_core_keymem_n371), .D(
        aes_core_keymem_n372), .Y(aes_core_round_key[22]) );
  AOI222X1 aes_core_keymem_U2477 ( .A0(aes_core_keymem_key_mem[310]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[54]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[182]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n231) );
  AOI222X1 aes_core_keymem_U2476 ( .A0(aes_core_keymem_key_mem[822]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[566]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[694]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n232) );
  AOI22X1 aes_core_keymem_U2475 ( .A0(aes_core_keymem_key_mem[1206]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1334]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n229) );
  NAND4X1 aes_core_keymem_U2474 ( .A(aes_core_keymem_n229), .B(
        aes_core_keymem_n230), .C(aes_core_keymem_n231), .D(
        aes_core_keymem_n232), .Y(aes_core_round_key[54]) );
  AOI222X1 aes_core_keymem_U2473 ( .A0(aes_core_keymem_key_mem[342]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[86]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[214]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n91) );
  AOI222X1 aes_core_keymem_U2472 ( .A0(aes_core_keymem_key_mem[854]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[598]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[726]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n92) );
  AOI22X1 aes_core_keymem_U2471 ( .A0(aes_core_keymem_key_mem[1238]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1366]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n89) );
  NAND4X1 aes_core_keymem_U2470 ( .A(aes_core_keymem_n89), .B(
        aes_core_keymem_n90), .C(aes_core_keymem_n91), .D(aes_core_keymem_n92), 
        .Y(aes_core_round_key[86]) );
  AOI222X1 aes_core_keymem_U2469 ( .A0(aes_core_keymem_key_mem[327]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[71]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[199]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n155) );
  AOI222X1 aes_core_keymem_U2468 ( .A0(aes_core_keymem_key_mem[839]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[583]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[711]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n156) );
  AOI22X1 aes_core_keymem_U2467 ( .A0(aes_core_keymem_key_mem[1223]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1351]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n153) );
  NAND4X1 aes_core_keymem_U2466 ( .A(aes_core_keymem_n153), .B(
        aes_core_keymem_n154), .C(aes_core_keymem_n155), .D(
        aes_core_keymem_n156), .Y(aes_core_round_key[71]) );
  AOI222X1 aes_core_keymem_U2464 ( .A0(aes_core_keymem_key_mem[311]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[55]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[183]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n227) );
  AOI222X1 aes_core_keymem_U2463 ( .A0(aes_core_keymem_key_mem[823]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[567]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[695]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n228) );
  AOI22X1 aes_core_keymem_U2462 ( .A0(aes_core_keymem_key_mem[1207]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1335]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n225) );
  NAND4X1 aes_core_keymem_U2461 ( .A(aes_core_keymem_n225), .B(
        aes_core_keymem_n226), .C(aes_core_keymem_n227), .D(
        aes_core_keymem_n228), .Y(aes_core_round_key[55]) );
  AOI222X1 aes_core_keymem_U2460 ( .A0(aes_core_keymem_key_mem[343]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[87]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[215]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n87) );
  AOI222X1 aes_core_keymem_U2459 ( .A0(aes_core_keymem_key_mem[855]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[599]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[727]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n88) );
  AOI22X1 aes_core_keymem_U2458 ( .A0(aes_core_keymem_key_mem[1239]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1367]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n85) );
  NAND4X1 aes_core_keymem_U2457 ( .A(aes_core_keymem_n85), .B(
        aes_core_keymem_n86), .C(aes_core_keymem_n87), .D(aes_core_keymem_n88), 
        .Y(aes_core_round_key[87]) );
  AOI222X1 aes_core_keymem_U2455 ( .A0(aes_core_keymem_key_mem[375]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[119]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[247]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n455) );
  AOI222X1 aes_core_keymem_U2453 ( .A0(aes_core_keymem_key_mem[887]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[631]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[759]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n456) );
  AOI22X1 aes_core_keymem_U2451 ( .A0(aes_core_keymem_key_mem[1271]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1399]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n453) );
  NAND4X1 aes_core_keymem_U2449 ( .A(aes_core_keymem_n453), .B(
        aes_core_keymem_n454), .C(aes_core_keymem_n455), .D(
        aes_core_keymem_n456), .Y(aes_core_round_key[119]) );
  AOI222X1 aes_core_keymem_U2447 ( .A0(aes_core_keymem_key_mem[279]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[23]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[151]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n367) );
  AOI222X1 aes_core_keymem_U2445 ( .A0(aes_core_keymem_key_mem[791]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[535]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[663]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n368) );
  AOI22X1 aes_core_keymem_U2443 ( .A0(aes_core_keymem_key_mem[1175]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1303]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n365) );
  NAND4X1 aes_core_keymem_U2442 ( .A(aes_core_keymem_n365), .B(
        aes_core_keymem_n366), .C(aes_core_keymem_n367), .D(
        aes_core_keymem_n368), .Y(aes_core_round_key[23]) );
  AOI222X1 aes_core_keymem_U2441 ( .A0(aes_core_keymem_key_mem[360]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[104]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[232]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n519) );
  AOI222X1 aes_core_keymem_U2440 ( .A0(aes_core_keymem_key_mem[872]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[616]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[744]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n520) );
  AOI22X1 aes_core_keymem_U2439 ( .A0(aes_core_keymem_key_mem[1256]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1384]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n517) );
  NAND4X1 aes_core_keymem_U2438 ( .A(aes_core_keymem_n517), .B(
        aes_core_keymem_n518), .C(aes_core_keymem_n519), .D(
        aes_core_keymem_n520), .Y(aes_core_round_key[104]) );
  AOI222X1 aes_core_keymem_U2437 ( .A0(aes_core_keymem_key_mem[296]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[40]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[168]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n291) );
  AOI222X1 aes_core_keymem_U2436 ( .A0(aes_core_keymem_key_mem[808]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[552]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[680]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n292) );
  AOI22X1 aes_core_keymem_U2435 ( .A0(aes_core_keymem_key_mem[1192]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1320]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n289) );
  NAND4X1 aes_core_keymem_U2434 ( .A(aes_core_keymem_n289), .B(
        aes_core_keymem_n290), .C(aes_core_keymem_n291), .D(
        aes_core_keymem_n292), .Y(aes_core_round_key[40]) );
  AOI222X1 aes_core_keymem_U2433 ( .A0(aes_core_keymem_key_mem[368]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[112]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[240]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n483) );
  AOI222X1 aes_core_keymem_U2432 ( .A0(aes_core_keymem_key_mem[880]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[624]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[752]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n484) );
  AOI22X1 aes_core_keymem_U2431 ( .A0(aes_core_keymem_key_mem[1264]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1392]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n481) );
  NAND4X1 aes_core_keymem_U2430 ( .A(aes_core_keymem_n481), .B(
        aes_core_keymem_n482), .C(aes_core_keymem_n483), .D(
        aes_core_keymem_n484), .Y(aes_core_round_key[112]) );
  AOI222X1 aes_core_keymem_U2429 ( .A0(aes_core_keymem_key_mem[272]), .A1(
        aes_core_keymem_n2719), .B0(aes_core_keymem_key_mem[16]), .B1(
        aes_core_keymem_n26), .C0(aes_core_keymem_key_mem[144]), .C1(
        aes_core_keymem_n2697), .Y(aes_core_keymem_n399) );
  AOI222X1 aes_core_keymem_U2428 ( .A0(aes_core_keymem_key_mem[784]), .A1(
        aes_core_keymem_n2752), .B0(aes_core_keymem_key_mem[528]), .B1(
        aes_core_keymem_n2741), .C0(aes_core_keymem_key_mem[656]), .C1(
        aes_core_keymem_n2730), .Y(aes_core_keymem_n400) );
  AOI22X1 aes_core_keymem_U2427 ( .A0(aes_core_keymem_key_mem[1168]), .A1(
        aes_core_keymem_n31), .B0(aes_core_keymem_key_mem[1296]), .B1(
        aes_core_keymem_n2644), .Y(aes_core_keymem_n397) );
  NAND4X1 aes_core_keymem_U2426 ( .A(aes_core_keymem_n397), .B(
        aes_core_keymem_n398), .C(aes_core_keymem_n399), .D(
        aes_core_keymem_n400), .Y(aes_core_round_key[16]) );
  AOI222X1 aes_core_keymem_U2425 ( .A0(aes_core_keymem_key_mem[304]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[48]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[176]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n259) );
  AOI222X1 aes_core_keymem_U2424 ( .A0(aes_core_keymem_key_mem[816]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[560]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[688]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n260) );
  AOI22X1 aes_core_keymem_U2423 ( .A0(aes_core_keymem_key_mem[1200]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1328]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n257) );
  NAND4X1 aes_core_keymem_U2422 ( .A(aes_core_keymem_n257), .B(
        aes_core_keymem_n258), .C(aes_core_keymem_n259), .D(
        aes_core_keymem_n260), .Y(aes_core_round_key[48]) );
  AOI222X1 aes_core_keymem_U2421 ( .A0(aes_core_keymem_key_mem[264]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[8]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[136]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n75) );
  AOI222X1 aes_core_keymem_U2420 ( .A0(aes_core_keymem_key_mem[776]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[520]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[648]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n76) );
  AOI22X1 aes_core_keymem_U2419 ( .A0(aes_core_keymem_key_mem[1160]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1288]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n73) );
  NAND4X1 aes_core_keymem_U2418 ( .A(aes_core_keymem_n73), .B(
        aes_core_keymem_n74), .C(aes_core_keymem_n75), .D(aes_core_keymem_n76), 
        .Y(aes_core_round_key[8]) );
  AOI222X1 aes_core_keymem_U2417 ( .A0(aes_core_keymem_key_mem[336]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[80]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[208]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n115) );
  AOI222X1 aes_core_keymem_U2416 ( .A0(aes_core_keymem_key_mem[848]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[592]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[720]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n116) );
  AOI22X1 aes_core_keymem_U2415 ( .A0(aes_core_keymem_key_mem[1232]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1360]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n113) );
  NAND4X1 aes_core_keymem_U2414 ( .A(aes_core_keymem_n113), .B(
        aes_core_keymem_n114), .C(aes_core_keymem_n115), .D(
        aes_core_keymem_n116), .Y(aes_core_round_key[80]) );
  AOI222X1 aes_core_keymem_U2413 ( .A0(aes_core_keymem_key_mem[305]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[49]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[177]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n255) );
  AOI222X1 aes_core_keymem_U2412 ( .A0(aes_core_keymem_key_mem[817]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[561]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[689]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n256) );
  AOI22X1 aes_core_keymem_U2411 ( .A0(aes_core_keymem_key_mem[1201]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1329]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n253) );
  NAND4X1 aes_core_keymem_U2410 ( .A(aes_core_keymem_n253), .B(
        aes_core_keymem_n254), .C(aes_core_keymem_n255), .D(
        aes_core_keymem_n256), .Y(aes_core_round_key[49]) );
  AOI222X1 aes_core_keymem_U2409 ( .A0(aes_core_keymem_key_mem[337]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[81]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[209]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n111) );
  AOI222X1 aes_core_keymem_U2408 ( .A0(aes_core_keymem_key_mem[849]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[593]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[721]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n112) );
  AOI22X1 aes_core_keymem_U2407 ( .A0(aes_core_keymem_key_mem[1233]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1361]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n109) );
  NAND4X1 aes_core_keymem_U2406 ( .A(aes_core_keymem_n109), .B(
        aes_core_keymem_n110), .C(aes_core_keymem_n111), .D(
        aes_core_keymem_n112), .Y(aes_core_round_key[81]) );
  AOI222X1 aes_core_keymem_U2405 ( .A0(aes_core_keymem_key_mem[369]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[113]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[241]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n479) );
  AOI222X1 aes_core_keymem_U2404 ( .A0(aes_core_keymem_key_mem[881]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[625]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[753]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n480) );
  AOI22X1 aes_core_keymem_U2403 ( .A0(aes_core_keymem_key_mem[1265]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1393]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n477) );
  NAND4X1 aes_core_keymem_U2402 ( .A(aes_core_keymem_n477), .B(
        aes_core_keymem_n478), .C(aes_core_keymem_n479), .D(
        aes_core_keymem_n480), .Y(aes_core_round_key[113]) );
  AOI222X1 aes_core_keymem_U2401 ( .A0(aes_core_keymem_key_mem[361]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[105]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[233]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n515) );
  AOI222X1 aes_core_keymem_U2400 ( .A0(aes_core_keymem_key_mem[873]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[617]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[745]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n516) );
  AOI22X1 aes_core_keymem_U2399 ( .A0(aes_core_keymem_key_mem[1257]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1385]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n513) );
  NAND4X1 aes_core_keymem_U2398 ( .A(aes_core_keymem_n513), .B(
        aes_core_keymem_n514), .C(aes_core_keymem_n515), .D(
        aes_core_keymem_n516), .Y(aes_core_round_key[105]) );
  AOI222X1 aes_core_keymem_U2397 ( .A0(aes_core_keymem_key_mem[329]), .A1(
        aes_core_keymem_n2724), .B0(aes_core_keymem_key_mem[73]), .B1(
        aes_core_keymem_n2713), .C0(aes_core_keymem_key_mem[201]), .C1(
        aes_core_keymem_n2702), .Y(aes_core_keymem_n147) );
  AOI222X1 aes_core_keymem_U2396 ( .A0(aes_core_keymem_key_mem[841]), .A1(
        aes_core_keymem_n2758), .B0(aes_core_keymem_key_mem[585]), .B1(
        aes_core_keymem_n2747), .C0(aes_core_keymem_key_mem[713]), .C1(
        aes_core_keymem_n2736), .Y(aes_core_keymem_n148) );
  AOI22X1 aes_core_keymem_U2395 ( .A0(aes_core_keymem_key_mem[1225]), .A1(
        aes_core_keymem_n2659), .B0(aes_core_keymem_key_mem[1353]), .B1(
        aes_core_keymem_n2649), .Y(aes_core_keymem_n145) );
  NAND4X1 aes_core_keymem_U2394 ( .A(aes_core_keymem_n145), .B(
        aes_core_keymem_n146), .C(aes_core_keymem_n147), .D(
        aes_core_keymem_n148), .Y(aes_core_round_key[73]) );
  AOI222X1 aes_core_keymem_U2393 ( .A0(aes_core_keymem_key_mem[273]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[17]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[145]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n395) );
  AOI222X1 aes_core_keymem_U2392 ( .A0(aes_core_keymem_key_mem[785]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[529]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[657]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n396) );
  AOI22X1 aes_core_keymem_U2391 ( .A0(aes_core_keymem_key_mem[1169]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1297]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n393) );
  NAND4X1 aes_core_keymem_U2390 ( .A(aes_core_keymem_n393), .B(
        aes_core_keymem_n394), .C(aes_core_keymem_n395), .D(
        aes_core_keymem_n396), .Y(aes_core_round_key[17]) );
  AOI222X1 aes_core_keymem_U2389 ( .A0(aes_core_keymem_key_mem[306]), .A1(
        aes_core_keymem_n2722), .B0(aes_core_keymem_key_mem[50]), .B1(
        aes_core_keymem_n2711), .C0(aes_core_keymem_key_mem[178]), .C1(
        aes_core_keymem_n2701), .Y(aes_core_keymem_n247) );
  AOI222X1 aes_core_keymem_U2388 ( .A0(aes_core_keymem_key_mem[818]), .A1(
        aes_core_keymem_n2756), .B0(aes_core_keymem_key_mem[562]), .B1(
        aes_core_keymem_n2745), .C0(aes_core_keymem_key_mem[690]), .C1(
        aes_core_keymem_n2734), .Y(aes_core_keymem_n248) );
  AOI22X1 aes_core_keymem_U2387 ( .A0(aes_core_keymem_key_mem[1202]), .A1(
        aes_core_keymem_n2657), .B0(aes_core_keymem_key_mem[1330]), .B1(
        aes_core_keymem_n2647), .Y(aes_core_keymem_n245) );
  NAND4X1 aes_core_keymem_U2386 ( .A(aes_core_keymem_n245), .B(
        aes_core_keymem_n246), .C(aes_core_keymem_n247), .D(
        aes_core_keymem_n248), .Y(aes_core_round_key[50]) );
  AOI222X1 aes_core_keymem_U2385 ( .A0(aes_core_keymem_key_mem[338]), .A1(
        aes_core_keymem_n2725), .B0(aes_core_keymem_key_mem[82]), .B1(
        aes_core_keymem_n2714), .C0(aes_core_keymem_key_mem[210]), .C1(
        aes_core_keymem_n2703), .Y(aes_core_keymem_n107) );
  AOI222X1 aes_core_keymem_U2384 ( .A0(aes_core_keymem_key_mem[850]), .A1(
        aes_core_keymem_n2759), .B0(aes_core_keymem_key_mem[594]), .B1(
        aes_core_keymem_n2748), .C0(aes_core_keymem_key_mem[722]), .C1(
        aes_core_keymem_n2737), .Y(aes_core_keymem_n108) );
  AOI22X1 aes_core_keymem_U2383 ( .A0(aes_core_keymem_key_mem[1234]), .A1(
        aes_core_keymem_n2660), .B0(aes_core_keymem_key_mem[1362]), .B1(
        aes_core_keymem_n2650), .Y(aes_core_keymem_n105) );
  NAND4X1 aes_core_keymem_U2382 ( .A(aes_core_keymem_n105), .B(
        aes_core_keymem_n106), .C(aes_core_keymem_n107), .D(
        aes_core_keymem_n108), .Y(aes_core_round_key[82]) );
  AOI222X1 aes_core_keymem_U2381 ( .A0(aes_core_keymem_key_mem[370]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[114]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[242]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n475) );
  AOI222X1 aes_core_keymem_U2380 ( .A0(aes_core_keymem_key_mem[882]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[626]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[754]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n476) );
  AOI22X1 aes_core_keymem_U2379 ( .A0(aes_core_keymem_key_mem[1266]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1394]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n473) );
  NAND4X1 aes_core_keymem_U2378 ( .A(aes_core_keymem_n473), .B(
        aes_core_keymem_n474), .C(aes_core_keymem_n475), .D(
        aes_core_keymem_n476), .Y(aes_core_round_key[114]) );
  AOI222X1 aes_core_keymem_U2377 ( .A0(aes_core_keymem_key_mem[274]), .A1(
        aes_core_keymem_n2720), .B0(aes_core_keymem_key_mem[18]), .B1(
        aes_core_keymem_n2708), .C0(aes_core_keymem_key_mem[146]), .C1(
        aes_core_keymem_n2698), .Y(aes_core_keymem_n391) );
  AOI222X1 aes_core_keymem_U2376 ( .A0(aes_core_keymem_key_mem[786]), .A1(
        aes_core_keymem_n2753), .B0(aes_core_keymem_key_mem[530]), .B1(
        aes_core_keymem_n2742), .C0(aes_core_keymem_key_mem[658]), .C1(
        aes_core_keymem_n2731), .Y(aes_core_keymem_n392) );
  AOI22X1 aes_core_keymem_U2375 ( .A0(aes_core_keymem_key_mem[1170]), .A1(
        aes_core_keymem_n2654), .B0(aes_core_keymem_key_mem[1298]), .B1(
        aes_core_keymem_n2645), .Y(aes_core_keymem_n389) );
  NAND4X1 aes_core_keymem_U2374 ( .A(aes_core_keymem_n389), .B(
        aes_core_keymem_n390), .C(aes_core_keymem_n391), .D(
        aes_core_keymem_n392), .Y(aes_core_round_key[18]) );
  AOI222X1 aes_core_keymem_U2373 ( .A0(aes_core_keymem_key_mem[371]), .A1(
        aes_core_keymem_n2718), .B0(aes_core_keymem_key_mem[115]), .B1(
        aes_core_keymem_n2707), .C0(aes_core_keymem_key_mem[243]), .C1(
        aes_core_keymem_n2696), .Y(aes_core_keymem_n471) );
  AOI222X1 aes_core_keymem_U2372 ( .A0(aes_core_keymem_key_mem[883]), .A1(
        aes_core_keymem_n2751), .B0(aes_core_keymem_key_mem[627]), .B1(
        aes_core_keymem_n2740), .C0(aes_core_keymem_key_mem[755]), .C1(
        aes_core_keymem_n2729), .Y(aes_core_keymem_n472) );
  AOI22X1 aes_core_keymem_U2371 ( .A0(aes_core_keymem_key_mem[1267]), .A1(
        aes_core_keymem_n2653), .B0(aes_core_keymem_key_mem[1395]), .B1(
        aes_core_keymem_n2643), .Y(aes_core_keymem_n469) );
  NAND4X1 aes_core_keymem_U2370 ( .A(aes_core_keymem_n469), .B(
        aes_core_keymem_n470), .C(aes_core_keymem_n471), .D(
        aes_core_keymem_n472), .Y(aes_core_round_key[115]) );
  AOI222X1 aes_core_keymem_U2369 ( .A0(aes_core_keymem_key_mem[290]), .A1(
        aes_core_keymem_n25), .B0(aes_core_keymem_key_mem[34]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[162]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n319) );
  AOI222X1 aes_core_keymem_U2368 ( .A0(aes_core_keymem_key_mem[802]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[546]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[674]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n320) );
  AOI22X1 aes_core_keymem_U2367 ( .A0(aes_core_keymem_key_mem[1186]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1314]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n317) );
  NAND4X1 aes_core_keymem_U2366 ( .A(aes_core_keymem_n317), .B(
        aes_core_keymem_n318), .C(aes_core_keymem_n319), .D(
        aes_core_keymem_n320), .Y(aes_core_round_key[34]) );
  AOI222X1 aes_core_keymem_U2365 ( .A0(aes_core_keymem_key_mem[259]), .A1(
        aes_core_keymem_n2721), .B0(aes_core_keymem_key_mem[3]), .B1(
        aes_core_keymem_n2710), .C0(aes_core_keymem_key_mem[131]), .C1(
        aes_core_keymem_n2700), .Y(aes_core_keymem_n295) );
  AOI222X1 aes_core_keymem_U2364 ( .A0(aes_core_keymem_key_mem[771]), .A1(
        aes_core_keymem_n2755), .B0(aes_core_keymem_key_mem[515]), .B1(
        aes_core_keymem_n2744), .C0(aes_core_keymem_key_mem[643]), .C1(
        aes_core_keymem_n2733), .Y(aes_core_keymem_n296) );
  AOI22X1 aes_core_keymem_U2363 ( .A0(aes_core_keymem_key_mem[1155]), .A1(
        aes_core_keymem_n2656), .B0(aes_core_keymem_key_mem[1283]), .B1(
        aes_core_keymem_n2646), .Y(aes_core_keymem_n293) );
  NAND4X1 aes_core_keymem_U2362 ( .A(aes_core_keymem_n293), .B(
        aes_core_keymem_n294), .C(aes_core_keymem_n295), .D(
        aes_core_keymem_n296), .Y(aes_core_round_key[3]) );
  AOI222X1 aes_core_keymem_U2361 ( .A0(aes_core_keymem_key_mem[289]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[33]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[161]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n323) );
  AOI222X1 aes_core_keymem_U2360 ( .A0(aes_core_keymem_key_mem[801]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[545]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[673]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n324) );
  AOI22X1 aes_core_keymem_U2359 ( .A0(aes_core_keymem_key_mem[1185]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1313]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n321) );
  NAND4X1 aes_core_keymem_U2358 ( .A(aes_core_keymem_n321), .B(
        aes_core_keymem_n322), .C(aes_core_keymem_n323), .D(
        aes_core_keymem_n324), .Y(aes_core_round_key[33]) );
  AOI222X1 aes_core_keymem_U2357 ( .A0(aes_core_keymem_key_mem[258]), .A1(
        aes_core_keymem_n2726), .B0(aes_core_keymem_key_mem[2]), .B1(
        aes_core_keymem_n2709), .C0(aes_core_keymem_key_mem[130]), .C1(
        aes_core_keymem_n2699), .Y(aes_core_keymem_n339) );
  AOI222X1 aes_core_keymem_U2356 ( .A0(aes_core_keymem_key_mem[770]), .A1(
        aes_core_keymem_n2754), .B0(aes_core_keymem_key_mem[514]), .B1(
        aes_core_keymem_n2743), .C0(aes_core_keymem_key_mem[642]), .C1(
        aes_core_keymem_n2732), .Y(aes_core_keymem_n340) );
  AOI22X1 aes_core_keymem_U2355 ( .A0(aes_core_keymem_key_mem[1154]), .A1(
        aes_core_keymem_n2655), .B0(aes_core_keymem_key_mem[1282]), .B1(
        aes_core_keymem_n32), .Y(aes_core_keymem_n337) );
  NAND4X1 aes_core_keymem_U2354 ( .A(aes_core_keymem_n337), .B(
        aes_core_keymem_n338), .C(aes_core_keymem_n339), .D(
        aes_core_keymem_n340), .Y(aes_core_round_key[2]) );
  AOI222X1 aes_core_keymem_U2353 ( .A0(aes_core_keymem_key_mem[266]), .A1(
        aes_core_keymem_n2717), .B0(aes_core_keymem_key_mem[10]), .B1(
        aes_core_keymem_n2706), .C0(aes_core_keymem_key_mem[138]), .C1(
        aes_core_keymem_n2695), .Y(aes_core_keymem_n495) );
  AOI222X1 aes_core_keymem_U2352 ( .A0(aes_core_keymem_key_mem[778]), .A1(
        aes_core_keymem_n2750), .B0(aes_core_keymem_key_mem[522]), .B1(
        aes_core_keymem_n2739), .C0(aes_core_keymem_key_mem[650]), .C1(
        aes_core_keymem_n2728), .Y(aes_core_keymem_n496) );
  AOI22X1 aes_core_keymem_U2351 ( .A0(aes_core_keymem_key_mem[1162]), .A1(
        aes_core_keymem_n2652), .B0(aes_core_keymem_key_mem[1290]), .B1(
        aes_core_keymem_n2642), .Y(aes_core_keymem_n493) );
  NAND4X1 aes_core_keymem_U2350 ( .A(aes_core_keymem_n493), .B(
        aes_core_keymem_n494), .C(aes_core_keymem_n495), .D(
        aes_core_keymem_n496), .Y(aes_core_round_key[10]) );
  INVX1 aes_core_keymem_U2349 ( .A(aes_core_enc_round_nr[1]), .Y(
        aes_core_keymem_n2772) );
  AND3X2 aes_core_keymem_U2348 ( .A(aes_core_enc_round_nr[0]), .B(
        aes_core_keymem_n2772), .C(aes_core_keymem_n542), .Y(
        aes_core_keymem_n31) );
  AOI222X1 aes_core_keymem_U2347 ( .A0(aes_core_keymem_key_mem[1120]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[480]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[992]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n46) );
  AOI222X1 aes_core_keymem_U2346 ( .A0(aes_core_keymem_key_mem[1121]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[481]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[993]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n42) );
  AOI222X1 aes_core_keymem_U2345 ( .A0(aes_core_keymem_key_mem[1033]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[393]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[905]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n19) );
  AOI222X1 aes_core_keymem_U2344 ( .A0(aes_core_keymem_key_mem[1123]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[483]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[995]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n34) );
  AOI222X1 aes_core_keymem_U2343 ( .A0(aes_core_keymem_key_mem[1122]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[482]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[994]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n38) );
  AOI222X1 aes_core_keymem_U2342 ( .A0(aes_core_keymem_key_mem[1119]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[479]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[991]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n50) );
  AOI222X1 aes_core_keymem_U2341 ( .A0(aes_core_keymem_key_mem[1117]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[477]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[989]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n58) );
  AOI222X1 aes_core_keymem_U2340 ( .A0(aes_core_keymem_key_mem[1118]), .A1(
        aes_core_keymem_n28), .B0(aes_core_keymem_key_mem[478]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[990]), .C1(
        aes_core_keymem_n2662), .Y(aes_core_keymem_n54) );
  AOI222X1 aes_core_keymem_U2339 ( .A0(aes_core_keymem_key_mem[1148]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[508]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[1020]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n430) );
  AOI222X1 aes_core_keymem_U2338 ( .A0(aes_core_keymem_key_mem[1052]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[412]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[924]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n346) );
  AOI222X1 aes_core_keymem_U2337 ( .A0(aes_core_keymem_key_mem[1084]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[444]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[956]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n202) );
  AOI222X1 aes_core_keymem_U2336 ( .A0(aes_core_keymem_key_mem[1116]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[476]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[988]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n62) );
  AOI222X1 aes_core_keymem_U2335 ( .A0(aes_core_keymem_key_mem[1113]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[473]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[985]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n78) );
  AOI222X1 aes_core_keymem_U2334 ( .A0(aes_core_keymem_key_mem[1145]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[505]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[1017]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n442) );
  AOI222X1 aes_core_keymem_U2333 ( .A0(aes_core_keymem_key_mem[1049]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[409]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[921]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n358) );
  AOI222X1 aes_core_keymem_U2332 ( .A0(aes_core_keymem_key_mem[1081]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[441]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[953]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n218) );
  AOI222X1 aes_core_keymem_U2331 ( .A0(aes_core_keymem_key_mem[1147]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[507]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[1019]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n434) );
  AOI222X1 aes_core_keymem_U2330 ( .A0(aes_core_keymem_key_mem[1051]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[411]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[923]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n350) );
  AOI222X1 aes_core_keymem_U2329 ( .A0(aes_core_keymem_key_mem[1115]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[475]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[987]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n66) );
  AOI222X1 aes_core_keymem_U2328 ( .A0(aes_core_keymem_key_mem[1083]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[443]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[955]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n210) );
  AOI222X1 aes_core_keymem_U2327 ( .A0(aes_core_keymem_key_mem[1089]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[449]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[961]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n182) );
  AOI222X1 aes_core_keymem_U2326 ( .A0(aes_core_keymem_key_mem[1066]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[426]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[938]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n282) );
  AOI222X1 aes_core_keymem_U2325 ( .A0(aes_core_keymem_key_mem[1131]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[491]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1003]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n506) );
  AOI222X1 aes_core_keymem_U2324 ( .A0(aes_core_keymem_key_mem[1059]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[419]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[931]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n314) );
  AOI222X1 aes_core_keymem_U2323 ( .A0(aes_core_keymem_key_mem[1028]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[388]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[900]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n250) );
  AOI222X1 aes_core_keymem_U2322 ( .A0(aes_core_keymem_key_mem[1133]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[493]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1005]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n498) );
  AOI222X1 aes_core_keymem_U2321 ( .A0(aes_core_keymem_key_mem[1061]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[421]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[933]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n306) );
  AOI222X1 aes_core_keymem_U2320 ( .A0(aes_core_keymem_key_mem[1029]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[389]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[901]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n206) );
  AOI222X1 aes_core_keymem_U2319 ( .A0(aes_core_keymem_key_mem[1134]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[494]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1006]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n490) );
  AOI222X1 aes_core_keymem_U2318 ( .A0(aes_core_keymem_key_mem[1062]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[422]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[934]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n302) );
  AOI222X1 aes_core_keymem_U2317 ( .A0(aes_core_keymem_key_mem[1030]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[390]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[902]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n162) );
  AOI222X1 aes_core_keymem_U2316 ( .A0(aes_core_keymem_key_mem[1135]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[495]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1007]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n486) );
  AOI222X1 aes_core_keymem_U2315 ( .A0(aes_core_keymem_key_mem[1063]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[423]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[935]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n298) );
  AOI222X1 aes_core_keymem_U2314 ( .A0(aes_core_keymem_key_mem[1024]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[384]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[896]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n538) );
  AOI222X1 aes_core_keymem_U2313 ( .A0(aes_core_keymem_key_mem[1090]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[450]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[962]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n178) );
  AOI222X1 aes_core_keymem_U2312 ( .A0(aes_core_keymem_key_mem[1067]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[427]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[939]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n278) );
  AOI222X1 aes_core_keymem_U2311 ( .A0(aes_core_keymem_key_mem[1132]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[492]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1004]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n502) );
  AOI222X1 aes_core_keymem_U2310 ( .A0(aes_core_keymem_key_mem[1060]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[420]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[932]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n310) );
  AOI222X1 aes_core_keymem_U2309 ( .A0(aes_core_keymem_key_mem[1036]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[396]), .B1(
        aes_core_keymem_n2682), .C0(aes_core_keymem_key_mem[908]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n414) );
  AOI222X1 aes_core_keymem_U2308 ( .A0(aes_core_keymem_key_mem[1092]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[452]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[964]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n170) );
  AOI222X1 aes_core_keymem_U2307 ( .A0(aes_core_keymem_key_mem[1069]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[429]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[941]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n270) );
  AOI222X1 aes_core_keymem_U2306 ( .A0(aes_core_keymem_key_mem[1125]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[485]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[997]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n530) );
  AOI222X1 aes_core_keymem_U2305 ( .A0(aes_core_keymem_key_mem[1093]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[453]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[965]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n166) );
  AOI222X1 aes_core_keymem_U2304 ( .A0(aes_core_keymem_key_mem[1070]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[430]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[942]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n266) );
  AOI222X1 aes_core_keymem_U2303 ( .A0(aes_core_keymem_key_mem[1126]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[486]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[998]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n526) );
  AOI222X1 aes_core_keymem_U2302 ( .A0(aes_core_keymem_key_mem[1094]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[454]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[966]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n158) );
  AOI222X1 aes_core_keymem_U2301 ( .A0(aes_core_keymem_key_mem[1071]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[431]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[943]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n262) );
  AOI222X1 aes_core_keymem_U2300 ( .A0(aes_core_keymem_key_mem[1127]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[487]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[999]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n522) );
  AOI222X1 aes_core_keymem_U2299 ( .A0(aes_core_keymem_key_mem[1088]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[448]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[960]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n186) );
  AOI222X1 aes_core_keymem_U2298 ( .A0(aes_core_keymem_key_mem[1065]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[425]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[937]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n286) );
  AOI222X1 aes_core_keymem_U2297 ( .A0(aes_core_keymem_key_mem[1130]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[490]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1002]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n510) );
  AOI222X1 aes_core_keymem_U2296 ( .A0(aes_core_keymem_key_mem[1075]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[435]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[947]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n242) );
  AOI222X1 aes_core_keymem_U2295 ( .A0(aes_core_keymem_key_mem[1108]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[468]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[980]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n98) );
  AOI222X1 aes_core_keymem_U2294 ( .A0(aes_core_keymem_key_mem[1124]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[484]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[996]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n534) );
  AOI222X1 aes_core_keymem_U2293 ( .A0(aes_core_keymem_key_mem[1100]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[460]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[972]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n134) );
  AOI222X1 aes_core_keymem_U2292 ( .A0(aes_core_keymem_key_mem[1037]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[397]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[909]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n410) );
  AOI222X1 aes_core_keymem_U2291 ( .A0(aes_core_keymem_key_mem[1102]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[462]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[974]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n126) );
  AOI222X1 aes_core_keymem_U2290 ( .A0(aes_core_keymem_key_mem[1039]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[399]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[911]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n402) );
  AOI222X1 aes_core_keymem_U2289 ( .A0(aes_core_keymem_key_mem[1096]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[456]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[968]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n150) );
  AOI222X1 aes_core_keymem_U2288 ( .A0(aes_core_keymem_key_mem[1098]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[458]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[970]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n142) );
  AOI222X1 aes_core_keymem_U2287 ( .A0(aes_core_keymem_key_mem[1035]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[395]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[907]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n450) );
  AOI222X1 aes_core_keymem_U2286 ( .A0(aes_core_keymem_key_mem[1091]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[451]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[963]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n174) );
  AOI222X1 aes_core_keymem_U2285 ( .A0(aes_core_keymem_key_mem[1068]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[428]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[940]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n274) );
  AOI222X1 aes_core_keymem_U2284 ( .A0(aes_core_keymem_key_mem[1141]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[501]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1013]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n462) );
  AOI222X1 aes_core_keymem_U2283 ( .A0(aes_core_keymem_key_mem[1038]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[398]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[910]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n406) );
  AOI222X1 aes_core_keymem_U2282 ( .A0(aes_core_keymem_key_mem[1103]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[463]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[975]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n122) );
  AOI222X1 aes_core_keymem_U2281 ( .A0(aes_core_keymem_key_mem[1031]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[391]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[903]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n118) );
  AOI222X1 aes_core_keymem_U2280 ( .A0(aes_core_keymem_key_mem[1107]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[467]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[979]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n102) );
  AOI222X1 aes_core_keymem_U2279 ( .A0(aes_core_keymem_key_mem[1140]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[500]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1012]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n466) );
  AOI222X1 aes_core_keymem_U2278 ( .A0(aes_core_keymem_key_mem[1044]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[404]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[916]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n378) );
  AOI222X1 aes_core_keymem_U2277 ( .A0(aes_core_keymem_key_mem[1056]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[416]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[928]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n326) );
  AOI222X1 aes_core_keymem_U2276 ( .A0(aes_core_keymem_key_mem[1025]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[385]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[897]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n382) );
  AOI222X1 aes_core_keymem_U2275 ( .A0(aes_core_keymem_key_mem[1099]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[459]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[971]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n138) );
  AOI222X1 aes_core_keymem_U2274 ( .A0(aes_core_keymem_key_mem[1043]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[403]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[915]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n386) );
  AOI222X1 aes_core_keymem_U2273 ( .A0(aes_core_keymem_key_mem[1076]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[436]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[948]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n238) );
  AOI222X1 aes_core_keymem_U2272 ( .A0(aes_core_keymem_key_mem[1101]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[461]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[973]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n130) );
  AOI222X1 aes_core_keymem_U2271 ( .A0(aes_core_keymem_key_mem[1045]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[405]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[917]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n374) );
  AOI222X1 aes_core_keymem_U2270 ( .A0(aes_core_keymem_key_mem[1077]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[437]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[949]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n234) );
  AOI222X1 aes_core_keymem_U2269 ( .A0(aes_core_keymem_key_mem[1109]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[469]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[981]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n94) );
  AOI222X1 aes_core_keymem_U2268 ( .A0(aes_core_keymem_key_mem[1142]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[502]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1014]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n458) );
  AOI222X1 aes_core_keymem_U2267 ( .A0(aes_core_keymem_key_mem[1046]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[406]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[918]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n370) );
  AOI222X1 aes_core_keymem_U2266 ( .A0(aes_core_keymem_key_mem[1078]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[438]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[950]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n230) );
  AOI222X1 aes_core_keymem_U2265 ( .A0(aes_core_keymem_key_mem[1110]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[470]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[982]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n90) );
  AOI222X1 aes_core_keymem_U2264 ( .A0(aes_core_keymem_key_mem[1095]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[455]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[967]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n154) );
  AOI222X1 aes_core_keymem_U2263 ( .A0(aes_core_keymem_key_mem[1079]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[439]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[951]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n226) );
  AOI222X1 aes_core_keymem_U2262 ( .A0(aes_core_keymem_key_mem[1111]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[471]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[983]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n86) );
  AOI222X1 aes_core_keymem_U2261 ( .A0(aes_core_keymem_key_mem[1143]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[503]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1015]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n454) );
  AOI222X1 aes_core_keymem_U2260 ( .A0(aes_core_keymem_key_mem[1047]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[407]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[919]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n366) );
  AOI222X1 aes_core_keymem_U2259 ( .A0(aes_core_keymem_key_mem[1128]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[488]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1000]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n518) );
  AOI222X1 aes_core_keymem_U2258 ( .A0(aes_core_keymem_key_mem[1064]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[424]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[936]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n290) );
  AOI222X1 aes_core_keymem_U2257 ( .A0(aes_core_keymem_key_mem[1136]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[496]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1008]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n482) );
  AOI222X1 aes_core_keymem_U2256 ( .A0(aes_core_keymem_key_mem[1040]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[400]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[912]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n398) );
  AOI222X1 aes_core_keymem_U2255 ( .A0(aes_core_keymem_key_mem[1072]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[432]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[944]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n258) );
  AOI222X1 aes_core_keymem_U2254 ( .A0(aes_core_keymem_key_mem[1032]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[392]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[904]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n74) );
  AOI222X1 aes_core_keymem_U2253 ( .A0(aes_core_keymem_key_mem[1104]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[464]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[976]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n114) );
  AOI222X1 aes_core_keymem_U2252 ( .A0(aes_core_keymem_key_mem[1073]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[433]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[945]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n254) );
  AOI222X1 aes_core_keymem_U2251 ( .A0(aes_core_keymem_key_mem[1105]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[465]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[977]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n110) );
  AOI222X1 aes_core_keymem_U2250 ( .A0(aes_core_keymem_key_mem[1137]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[497]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1009]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n478) );
  AOI222X1 aes_core_keymem_U2249 ( .A0(aes_core_keymem_key_mem[1129]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[489]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[1001]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n514) );
  AOI222X1 aes_core_keymem_U2248 ( .A0(aes_core_keymem_key_mem[1097]), .A1(
        aes_core_keymem_n2692), .B0(aes_core_keymem_key_mem[457]), .B1(
        aes_core_keymem_n2680), .C0(aes_core_keymem_key_mem[969]), .C1(
        aes_core_keymem_n2671), .Y(aes_core_keymem_n146) );
  AOI222X1 aes_core_keymem_U2247 ( .A0(aes_core_keymem_key_mem[1041]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[401]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[913]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n394) );
  AOI222X1 aes_core_keymem_U2246 ( .A0(aes_core_keymem_key_mem[1074]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[434]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[946]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n246) );
  AOI222X1 aes_core_keymem_U2245 ( .A0(aes_core_keymem_key_mem[1106]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[466]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[978]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n106) );
  AOI222X1 aes_core_keymem_U2244 ( .A0(aes_core_keymem_key_mem[1138]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[498]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1010]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n474) );
  AOI222X1 aes_core_keymem_U2243 ( .A0(aes_core_keymem_key_mem[1042]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[402]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[914]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n390) );
  AOI222X1 aes_core_keymem_U2242 ( .A0(aes_core_keymem_key_mem[1139]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[499]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1011]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n470) );
  AOI222X1 aes_core_keymem_U2241 ( .A0(aes_core_keymem_key_mem[1058]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[418]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[930]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n318) );
  AOI222X1 aes_core_keymem_U2240 ( .A0(aes_core_keymem_key_mem[1027]), .A1(
        aes_core_keymem_n2689), .B0(aes_core_keymem_key_mem[387]), .B1(
        aes_core_keymem_n2677), .C0(aes_core_keymem_key_mem[899]), .C1(
        aes_core_keymem_n2668), .Y(aes_core_keymem_n294) );
  AOI222X1 aes_core_keymem_U2239 ( .A0(aes_core_keymem_key_mem[1057]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[417]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[929]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n322) );
  AOI222X1 aes_core_keymem_U2238 ( .A0(aes_core_keymem_key_mem[1026]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[386]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[898]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n338) );
  AOI222X1 aes_core_keymem_U2237 ( .A0(aes_core_keymem_key_mem[1034]), .A1(
        aes_core_keymem_n2684), .B0(aes_core_keymem_key_mem[394]), .B1(
        aes_core_keymem_n2673), .C0(aes_core_keymem_key_mem[906]), .C1(
        aes_core_keymem_n2663), .Y(aes_core_keymem_n494) );
  AOI222X1 aes_core_keymem_U2236 ( .A0(aes_core_keymem_key_mem[1053]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[413]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[925]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n342) );
  AOI222X1 aes_core_keymem_U2235 ( .A0(aes_core_keymem_key_mem[1054]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[414]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[926]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n334) );
  AOI222X1 aes_core_keymem_U2234 ( .A0(aes_core_keymem_key_mem[1055]), .A1(
        aes_core_keymem_n2688), .B0(aes_core_keymem_key_mem[415]), .B1(
        aes_core_keymem_n2676), .C0(aes_core_keymem_key_mem[927]), .C1(
        aes_core_keymem_n2667), .Y(aes_core_keymem_n330) );
  AOI222X1 aes_core_keymem_U2233 ( .A0(aes_core_keymem_key_mem[1085]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[445]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[957]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n198) );
  AOI222X1 aes_core_keymem_U2232 ( .A0(aes_core_keymem_key_mem[1086]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[446]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[958]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n194) );
  AOI222X1 aes_core_keymem_U2231 ( .A0(aes_core_keymem_key_mem[1087]), .A1(
        aes_core_keymem_n2691), .B0(aes_core_keymem_key_mem[447]), .B1(
        aes_core_keymem_n2679), .C0(aes_core_keymem_key_mem[959]), .C1(
        aes_core_keymem_n2670), .Y(aes_core_keymem_n190) );
  AOI222X1 aes_core_keymem_U2230 ( .A0(aes_core_keymem_key_mem[1080]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[440]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[952]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n222) );
  AOI222X1 aes_core_keymem_U2229 ( .A0(aes_core_keymem_key_mem[1149]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[509]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[1021]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n426) );
  AOI222X1 aes_core_keymem_U2228 ( .A0(aes_core_keymem_key_mem[1150]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[510]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[1022]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n422) );
  AOI222X1 aes_core_keymem_U2227 ( .A0(aes_core_keymem_key_mem[1151]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[511]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[1023]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n418) );
  AOI222X1 aes_core_keymem_U2226 ( .A0(aes_core_keymem_key_mem[1144]), .A1(
        aes_core_keymem_n2685), .B0(aes_core_keymem_key_mem[504]), .B1(
        aes_core_keymem_n2674), .C0(aes_core_keymem_key_mem[1016]), .C1(
        aes_core_keymem_n2664), .Y(aes_core_keymem_n446) );
  AOI222X1 aes_core_keymem_U2225 ( .A0(aes_core_keymem_key_mem[1048]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[408]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[920]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n362) );
  AOI222X1 aes_core_keymem_U2224 ( .A0(aes_core_keymem_key_mem[1112]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[472]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[984]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n82) );
  AOI222X1 aes_core_keymem_U2223 ( .A0(aes_core_keymem_key_mem[1082]), .A1(
        aes_core_keymem_n2690), .B0(aes_core_keymem_key_mem[442]), .B1(
        aes_core_keymem_n2678), .C0(aes_core_keymem_key_mem[954]), .C1(
        aes_core_keymem_n2669), .Y(aes_core_keymem_n214) );
  AOI222X1 aes_core_keymem_U2222 ( .A0(aes_core_keymem_key_mem[1114]), .A1(
        aes_core_keymem_n2693), .B0(aes_core_keymem_key_mem[474]), .B1(
        aes_core_keymem_n2681), .C0(aes_core_keymem_key_mem[986]), .C1(
        aes_core_keymem_n2672), .Y(aes_core_keymem_n70) );
  AOI222X1 aes_core_keymem_U2221 ( .A0(aes_core_keymem_key_mem[1146]), .A1(
        aes_core_keymem_n2686), .B0(aes_core_keymem_key_mem[506]), .B1(
        aes_core_keymem_n29), .C0(aes_core_keymem_key_mem[1018]), .C1(
        aes_core_keymem_n2665), .Y(aes_core_keymem_n438) );
  AOI222X1 aes_core_keymem_U2220 ( .A0(aes_core_keymem_key_mem[1050]), .A1(
        aes_core_keymem_n2687), .B0(aes_core_keymem_key_mem[410]), .B1(
        aes_core_keymem_n2675), .C0(aes_core_keymem_key_mem[922]), .C1(
        aes_core_keymem_n2666), .Y(aes_core_keymem_n354) );
  OAI2BB2X1 aes_core_keymem_U2219 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1011]), .Y(aes_core_keymem_n993) );
  OAI2BB2X1 aes_core_keymem_U2218 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1139]), .Y(aes_core_keymem_n994) );
  OAI2BB2X1 aes_core_keymem_U2217 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1267]), .Y(aes_core_keymem_n995) );
  OAI2BB2X1 aes_core_keymem_U2216 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1395]), .Y(aes_core_keymem_n996) );
  OAI2BB2X1 aes_core_keymem_U2215 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1010]), .Y(aes_core_keymem_n1005) );
  OAI2BB2X1 aes_core_keymem_U2214 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1138]), .Y(aes_core_keymem_n1006) );
  OAI2BB2X1 aes_core_keymem_U2213 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1266]), .Y(aes_core_keymem_n1007) );
  OAI2BB2X1 aes_core_keymem_U2212 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1394]), .Y(aes_core_keymem_n1008) );
  OAI2BB2X1 aes_core_keymem_U2211 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1008]), .Y(aes_core_keymem_n1029) );
  OAI2BB2X1 aes_core_keymem_U2210 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1136]), .Y(aes_core_keymem_n1030) );
  OAI2BB2X1 aes_core_keymem_U2209 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1264]), .Y(aes_core_keymem_n1031) );
  OAI2BB2X1 aes_core_keymem_U2208 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1392]), .Y(aes_core_keymem_n1032) );
  OAI2BB2X1 aes_core_keymem_U2207 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[997]), .Y(aes_core_keymem_n1161) );
  OAI2BB2X1 aes_core_keymem_U2206 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1125]), .Y(aes_core_keymem_n1162) );
  OAI2BB2X1 aes_core_keymem_U2205 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1253]), .Y(aes_core_keymem_n1163) );
  OAI2BB2X1 aes_core_keymem_U2204 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1381]), .Y(aes_core_keymem_n1164) );
  OAI2BB2X1 aes_core_keymem_U2203 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[993]), .Y(aes_core_keymem_n1209) );
  OAI2BB2X1 aes_core_keymem_U2202 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1121]), .Y(aes_core_keymem_n1210) );
  OAI2BB2X1 aes_core_keymem_U2201 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1249]), .Y(aes_core_keymem_n1211) );
  OAI2BB2X1 aes_core_keymem_U2200 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1377]), .Y(aes_core_keymem_n1212) );
  OAI2BB2X1 aes_core_keymem_U2199 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1023]), .Y(aes_core_keymem_n849) );
  OAI2BB2X1 aes_core_keymem_U2198 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1151]), .Y(aes_core_keymem_n850) );
  OAI2BB2X1 aes_core_keymem_U2197 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1279]), .Y(aes_core_keymem_n851) );
  OAI2BB2X1 aes_core_keymem_U2196 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1407]), .Y(aes_core_keymem_n852) );
  OAI2BB2X1 aes_core_keymem_U2195 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1022]), .Y(aes_core_keymem_n861) );
  OAI2BB2X1 aes_core_keymem_U2194 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1150]), .Y(aes_core_keymem_n862) );
  OAI2BB2X1 aes_core_keymem_U2193 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1278]), .Y(aes_core_keymem_n863) );
  OAI2BB2X1 aes_core_keymem_U2192 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1406]), .Y(aes_core_keymem_n864) );
  OAI2BB2X1 aes_core_keymem_U2191 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1021]), .Y(aes_core_keymem_n873) );
  OAI2BB2X1 aes_core_keymem_U2190 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1149]), .Y(aes_core_keymem_n874) );
  OAI2BB2X1 aes_core_keymem_U2189 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1277]), .Y(aes_core_keymem_n875) );
  OAI2BB2X1 aes_core_keymem_U2188 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1405]), .Y(aes_core_keymem_n876) );
  OAI2BB2X1 aes_core_keymem_U2187 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1020]), .Y(aes_core_keymem_n885) );
  OAI2BB2X1 aes_core_keymem_U2186 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1148]), .Y(aes_core_keymem_n886) );
  OAI2BB2X1 aes_core_keymem_U2185 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1276]), .Y(aes_core_keymem_n887) );
  OAI2BB2X1 aes_core_keymem_U2184 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1404]), .Y(aes_core_keymem_n888) );
  OAI2BB2X1 aes_core_keymem_U2183 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1019]), .Y(aes_core_keymem_n897) );
  OAI2BB2X1 aes_core_keymem_U2182 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1147]), .Y(aes_core_keymem_n898) );
  OAI2BB2X1 aes_core_keymem_U2181 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1275]), .Y(aes_core_keymem_n899) );
  OAI2BB2X1 aes_core_keymem_U2180 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1403]), .Y(aes_core_keymem_n900) );
  OAI2BB2X1 aes_core_keymem_U2179 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[1018]), .Y(aes_core_keymem_n909) );
  OAI2BB2X1 aes_core_keymem_U2178 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1146]), .Y(aes_core_keymem_n910) );
  OAI2BB2X1 aes_core_keymem_U2177 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1274]), .Y(aes_core_keymem_n911) );
  OAI2BB2X1 aes_core_keymem_U2176 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1402]), .Y(aes_core_keymem_n912) );
  OAI2BB2X1 aes_core_keymem_U2175 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[1017]), .Y(aes_core_keymem_n921) );
  OAI2BB2X1 aes_core_keymem_U2174 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1145]), .Y(aes_core_keymem_n922) );
  OAI2BB2X1 aes_core_keymem_U2173 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1273]), .Y(aes_core_keymem_n923) );
  OAI2BB2X1 aes_core_keymem_U2172 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1401]), .Y(aes_core_keymem_n924) );
  OAI2BB2X1 aes_core_keymem_U2171 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1016]), .Y(aes_core_keymem_n933) );
  OAI2BB2X1 aes_core_keymem_U2170 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1144]), .Y(aes_core_keymem_n934) );
  OAI2BB2X1 aes_core_keymem_U2169 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1272]), .Y(aes_core_keymem_n935) );
  OAI2BB2X1 aes_core_keymem_U2168 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1400]), .Y(aes_core_keymem_n936) );
  OAI2BB2X1 aes_core_keymem_U2167 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1015]), .Y(aes_core_keymem_n945) );
  OAI2BB2X1 aes_core_keymem_U2166 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1143]), .Y(aes_core_keymem_n946) );
  OAI2BB2X1 aes_core_keymem_U2165 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1271]), .Y(aes_core_keymem_n947) );
  OAI2BB2X1 aes_core_keymem_U2164 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1399]), .Y(aes_core_keymem_n948) );
  OAI2BB2X1 aes_core_keymem_U2163 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1014]), .Y(aes_core_keymem_n957) );
  OAI2BB2X1 aes_core_keymem_U2162 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1142]), .Y(aes_core_keymem_n958) );
  OAI2BB2X1 aes_core_keymem_U2161 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1270]), .Y(aes_core_keymem_n959) );
  OAI2BB2X1 aes_core_keymem_U2160 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1398]), .Y(aes_core_keymem_n960) );
  OAI2BB2X1 aes_core_keymem_U2159 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1013]), .Y(aes_core_keymem_n969) );
  OAI2BB2X1 aes_core_keymem_U2158 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1141]), .Y(aes_core_keymem_n970) );
  OAI2BB2X1 aes_core_keymem_U2157 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1269]), .Y(aes_core_keymem_n971) );
  OAI2BB2X1 aes_core_keymem_U2156 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1397]), .Y(aes_core_keymem_n972) );
  OAI2BB2X1 aes_core_keymem_U2155 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n2626), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1012]), .Y(aes_core_keymem_n981) );
  OAI2BB2X1 aes_core_keymem_U2154 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n2610), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1140]), .Y(aes_core_keymem_n982) );
  OAI2BB2X1 aes_core_keymem_U2153 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n2593), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1268]), .Y(aes_core_keymem_n983) );
  OAI2BB2X1 aes_core_keymem_U2152 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n2506), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1396]), .Y(aes_core_keymem_n984) );
  OAI2BB2X1 aes_core_keymem_U2151 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1009]), .Y(aes_core_keymem_n1017) );
  OAI2BB2X1 aes_core_keymem_U2150 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1137]), .Y(aes_core_keymem_n1018) );
  OAI2BB2X1 aes_core_keymem_U2149 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1265]), .Y(aes_core_keymem_n1019) );
  OAI2BB2X1 aes_core_keymem_U2148 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1393]), .Y(aes_core_keymem_n1020) );
  OAI2BB2X1 aes_core_keymem_U2147 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1007]), .Y(aes_core_keymem_n1041) );
  OAI2BB2X1 aes_core_keymem_U2146 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1135]), .Y(aes_core_keymem_n1042) );
  OAI2BB2X1 aes_core_keymem_U2145 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1263]), .Y(aes_core_keymem_n1043) );
  OAI2BB2X1 aes_core_keymem_U2144 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1391]), .Y(aes_core_keymem_n1044) );
  OAI2BB2X1 aes_core_keymem_U2143 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[1006]), .Y(aes_core_keymem_n1053) );
  OAI2BB2X1 aes_core_keymem_U2142 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1134]), .Y(aes_core_keymem_n1054) );
  OAI2BB2X1 aes_core_keymem_U2141 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1262]), .Y(aes_core_keymem_n1055) );
  OAI2BB2X1 aes_core_keymem_U2140 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1390]), .Y(aes_core_keymem_n1056) );
  OAI2BB2X1 aes_core_keymem_U2139 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1005]), .Y(aes_core_keymem_n1065) );
  OAI2BB2X1 aes_core_keymem_U2138 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1133]), .Y(aes_core_keymem_n1066) );
  OAI2BB2X1 aes_core_keymem_U2137 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1261]), .Y(aes_core_keymem_n1067) );
  OAI2BB2X1 aes_core_keymem_U2136 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1389]), .Y(aes_core_keymem_n1068) );
  OAI2BB2X1 aes_core_keymem_U2135 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1004]), .Y(aes_core_keymem_n1077) );
  OAI2BB2X1 aes_core_keymem_U2134 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1132]), .Y(aes_core_keymem_n1078) );
  OAI2BB2X1 aes_core_keymem_U2133 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1260]), .Y(aes_core_keymem_n1079) );
  OAI2BB2X1 aes_core_keymem_U2132 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1388]), .Y(aes_core_keymem_n1080) );
  OAI2BB2X1 aes_core_keymem_U2131 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1003]), .Y(aes_core_keymem_n1089) );
  OAI2BB2X1 aes_core_keymem_U2130 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1131]), .Y(aes_core_keymem_n1090) );
  OAI2BB2X1 aes_core_keymem_U2129 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1259]), .Y(aes_core_keymem_n1091) );
  OAI2BB2X1 aes_core_keymem_U2128 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1387]), .Y(aes_core_keymem_n1092) );
  OAI2BB2X1 aes_core_keymem_U2127 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1002]), .Y(aes_core_keymem_n1101) );
  OAI2BB2X1 aes_core_keymem_U2126 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1130]), .Y(aes_core_keymem_n1102) );
  OAI2BB2X1 aes_core_keymem_U2125 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1258]), .Y(aes_core_keymem_n1103) );
  OAI2BB2X1 aes_core_keymem_U2124 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1386]), .Y(aes_core_keymem_n1104) );
  OAI2BB2X1 aes_core_keymem_U2123 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1001]), .Y(aes_core_keymem_n1113) );
  OAI2BB2X1 aes_core_keymem_U2122 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1129]), .Y(aes_core_keymem_n1114) );
  OAI2BB2X1 aes_core_keymem_U2121 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1257]), .Y(aes_core_keymem_n1115) );
  OAI2BB2X1 aes_core_keymem_U2120 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1385]), .Y(aes_core_keymem_n1116) );
  OAI2BB2X1 aes_core_keymem_U2119 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[1000]), .Y(aes_core_keymem_n1125) );
  OAI2BB2X1 aes_core_keymem_U2118 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1128]), .Y(aes_core_keymem_n1126) );
  OAI2BB2X1 aes_core_keymem_U2117 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1256]), .Y(aes_core_keymem_n1127) );
  OAI2BB2X1 aes_core_keymem_U2116 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1384]), .Y(aes_core_keymem_n1128) );
  OAI2BB2X1 aes_core_keymem_U2115 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n2627), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[999]), .Y(aes_core_keymem_n1137) );
  OAI2BB2X1 aes_core_keymem_U2114 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n2611), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1127]), .Y(aes_core_keymem_n1138) );
  OAI2BB2X1 aes_core_keymem_U2113 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n2594), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1255]), .Y(aes_core_keymem_n1139) );
  OAI2BB2X1 aes_core_keymem_U2112 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n2507), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1383]), .Y(aes_core_keymem_n1140) );
  OAI2BB2X1 aes_core_keymem_U2111 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[998]), .Y(aes_core_keymem_n1149) );
  OAI2BB2X1 aes_core_keymem_U2110 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1126]), .Y(aes_core_keymem_n1150) );
  OAI2BB2X1 aes_core_keymem_U2109 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1254]), .Y(aes_core_keymem_n1151) );
  OAI2BB2X1 aes_core_keymem_U2108 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1382]), .Y(aes_core_keymem_n1152) );
  OAI2BB2X1 aes_core_keymem_U2107 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[996]), .Y(aes_core_keymem_n1173) );
  OAI2BB2X1 aes_core_keymem_U2106 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1124]), .Y(aes_core_keymem_n1174) );
  OAI2BB2X1 aes_core_keymem_U2105 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1252]), .Y(aes_core_keymem_n1175) );
  OAI2BB2X1 aes_core_keymem_U2104 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1380]), .Y(aes_core_keymem_n1176) );
  OAI2BB2X1 aes_core_keymem_U2103 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[995]), .Y(aes_core_keymem_n1185) );
  OAI2BB2X1 aes_core_keymem_U2102 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1123]), .Y(aes_core_keymem_n1186) );
  OAI2BB2X1 aes_core_keymem_U2101 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1251]), .Y(aes_core_keymem_n1187) );
  OAI2BB2X1 aes_core_keymem_U2100 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1379]), .Y(aes_core_keymem_n1188) );
  OAI2BB2X1 aes_core_keymem_U2099 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[994]), .Y(aes_core_keymem_n1197) );
  OAI2BB2X1 aes_core_keymem_U2098 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1122]), .Y(aes_core_keymem_n1198) );
  OAI2BB2X1 aes_core_keymem_U2097 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1250]), .Y(aes_core_keymem_n1199) );
  OAI2BB2X1 aes_core_keymem_U2096 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1378]), .Y(aes_core_keymem_n1200) );
  OAI2BB2X1 aes_core_keymem_U2095 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[992]), .Y(aes_core_keymem_n1221) );
  OAI2BB2X1 aes_core_keymem_U2094 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1120]), .Y(aes_core_keymem_n1222) );
  OAI2BB2X1 aes_core_keymem_U2093 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1248]), .Y(aes_core_keymem_n1223) );
  OAI2BB2X1 aes_core_keymem_U2092 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1376]), .Y(aes_core_keymem_n1224) );
  OAI2BB2X1 aes_core_keymem_U2091 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[990]), .Y(aes_core_keymem_n1245) );
  OAI2BB2X1 aes_core_keymem_U2090 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1118]), .Y(aes_core_keymem_n1246) );
  OAI2BB2X1 aes_core_keymem_U2089 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1246]), .Y(aes_core_keymem_n1247) );
  OAI2BB2X1 aes_core_keymem_U2088 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1374]), .Y(aes_core_keymem_n1248) );
  OAI2BB2X1 aes_core_keymem_U2087 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[989]), .Y(aes_core_keymem_n1257) );
  OAI2BB2X1 aes_core_keymem_U2086 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1117]), .Y(aes_core_keymem_n1258) );
  OAI2BB2X1 aes_core_keymem_U2085 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1245]), .Y(aes_core_keymem_n1259) );
  OAI2BB2X1 aes_core_keymem_U2084 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1373]), .Y(aes_core_keymem_n1260) );
  OAI2BB2X1 aes_core_keymem_U2083 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[988]), .Y(aes_core_keymem_n1269) );
  OAI2BB2X1 aes_core_keymem_U2082 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1116]), .Y(aes_core_keymem_n1270) );
  OAI2BB2X1 aes_core_keymem_U2081 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1244]), .Y(aes_core_keymem_n1271) );
  OAI2BB2X1 aes_core_keymem_U2080 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1372]), .Y(aes_core_keymem_n1272) );
  OAI2BB2X1 aes_core_keymem_U2079 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[987]), .Y(aes_core_keymem_n1281) );
  OAI2BB2X1 aes_core_keymem_U2078 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1115]), .Y(aes_core_keymem_n1282) );
  OAI2BB2X1 aes_core_keymem_U2077 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1243]), .Y(aes_core_keymem_n1283) );
  OAI2BB2X1 aes_core_keymem_U2076 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1371]), .Y(aes_core_keymem_n1284) );
  OAI2BB2X1 aes_core_keymem_U2075 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[986]), .Y(aes_core_keymem_n1293) );
  OAI2BB2X1 aes_core_keymem_U2074 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1114]), .Y(aes_core_keymem_n1294) );
  OAI2BB2X1 aes_core_keymem_U2073 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1242]), .Y(aes_core_keymem_n1295) );
  OAI2BB2X1 aes_core_keymem_U2072 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1370]), .Y(aes_core_keymem_n1296) );
  OAI2BB2X1 aes_core_keymem_U2071 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[985]), .Y(aes_core_keymem_n1305) );
  OAI2BB2X1 aes_core_keymem_U2070 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1113]), .Y(aes_core_keymem_n1306) );
  OAI2BB2X1 aes_core_keymem_U2069 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1241]), .Y(aes_core_keymem_n1307) );
  OAI2BB2X1 aes_core_keymem_U2068 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1369]), .Y(aes_core_keymem_n1308) );
  OAI2BB2X1 aes_core_keymem_U2067 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[984]), .Y(aes_core_keymem_n1317) );
  OAI2BB2X1 aes_core_keymem_U2066 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1112]), .Y(aes_core_keymem_n1318) );
  OAI2BB2X1 aes_core_keymem_U2065 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1240]), .Y(aes_core_keymem_n1319) );
  OAI2BB2X1 aes_core_keymem_U2064 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1368]), .Y(aes_core_keymem_n1320) );
  OAI2BB2X1 aes_core_keymem_U2063 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[983]), .Y(aes_core_keymem_n1329) );
  OAI2BB2X1 aes_core_keymem_U2062 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1111]), .Y(aes_core_keymem_n1330) );
  OAI2BB2X1 aes_core_keymem_U2061 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1239]), .Y(aes_core_keymem_n1331) );
  OAI2BB2X1 aes_core_keymem_U2060 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1367]), .Y(aes_core_keymem_n1332) );
  OAI2BB2X1 aes_core_keymem_U2059 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[982]), .Y(aes_core_keymem_n1341) );
  OAI2BB2X1 aes_core_keymem_U2058 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1110]), .Y(aes_core_keymem_n1342) );
  OAI2BB2X1 aes_core_keymem_U2057 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1238]), .Y(aes_core_keymem_n1343) );
  OAI2BB2X1 aes_core_keymem_U2056 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1366]), .Y(aes_core_keymem_n1344) );
  OAI2BB2X1 aes_core_keymem_U2055 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[981]), .Y(aes_core_keymem_n1353) );
  OAI2BB2X1 aes_core_keymem_U2054 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1109]), .Y(aes_core_keymem_n1354) );
  OAI2BB2X1 aes_core_keymem_U2053 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1237]), .Y(aes_core_keymem_n1355) );
  OAI2BB2X1 aes_core_keymem_U2052 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1365]), .Y(aes_core_keymem_n1356) );
  OAI2BB2X1 aes_core_keymem_U2051 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[980]), .Y(aes_core_keymem_n1365) );
  OAI2BB2X1 aes_core_keymem_U2050 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1108]), .Y(aes_core_keymem_n1366) );
  OAI2BB2X1 aes_core_keymem_U2049 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1236]), .Y(aes_core_keymem_n1367) );
  OAI2BB2X1 aes_core_keymem_U2048 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1364]), .Y(aes_core_keymem_n1368) );
  OAI2BB2X1 aes_core_keymem_U2047 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[979]), .Y(aes_core_keymem_n1377) );
  OAI2BB2X1 aes_core_keymem_U2046 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1107]), .Y(aes_core_keymem_n1378) );
  OAI2BB2X1 aes_core_keymem_U2045 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1235]), .Y(aes_core_keymem_n1379) );
  OAI2BB2X1 aes_core_keymem_U2044 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1363]), .Y(aes_core_keymem_n1380) );
  OAI2BB2X1 aes_core_keymem_U2043 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[978]), .Y(aes_core_keymem_n1389) );
  OAI2BB2X1 aes_core_keymem_U2042 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1106]), .Y(aes_core_keymem_n1390) );
  OAI2BB2X1 aes_core_keymem_U2041 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1234]), .Y(aes_core_keymem_n1391) );
  OAI2BB2X1 aes_core_keymem_U2040 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1362]), .Y(aes_core_keymem_n1392) );
  OAI2BB2X1 aes_core_keymem_U2039 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[977]), .Y(aes_core_keymem_n1401) );
  OAI2BB2X1 aes_core_keymem_U2038 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1105]), .Y(aes_core_keymem_n1402) );
  OAI2BB2X1 aes_core_keymem_U2037 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1233]), .Y(aes_core_keymem_n1403) );
  OAI2BB2X1 aes_core_keymem_U2036 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1361]), .Y(aes_core_keymem_n1404) );
  OAI2BB2X1 aes_core_keymem_U2035 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[976]), .Y(aes_core_keymem_n1413) );
  OAI2BB2X1 aes_core_keymem_U2034 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1104]), .Y(aes_core_keymem_n1414) );
  OAI2BB2X1 aes_core_keymem_U2033 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1232]), .Y(aes_core_keymem_n1415) );
  OAI2BB2X1 aes_core_keymem_U2032 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1360]), .Y(aes_core_keymem_n1416) );
  OAI2BB2X1 aes_core_keymem_U2031 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[974]), .Y(aes_core_keymem_n1437) );
  OAI2BB2X1 aes_core_keymem_U2030 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1102]), .Y(aes_core_keymem_n1438) );
  OAI2BB2X1 aes_core_keymem_U2029 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1230]), .Y(aes_core_keymem_n1439) );
  OAI2BB2X1 aes_core_keymem_U2028 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1358]), .Y(aes_core_keymem_n1440) );
  OAI2BB2X1 aes_core_keymem_U2027 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[973]), .Y(aes_core_keymem_n1449) );
  OAI2BB2X1 aes_core_keymem_U2026 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1101]), .Y(aes_core_keymem_n1450) );
  OAI2BB2X1 aes_core_keymem_U2025 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1229]), .Y(aes_core_keymem_n1451) );
  OAI2BB2X1 aes_core_keymem_U2024 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1357]), .Y(aes_core_keymem_n1452) );
  OAI2BB2X1 aes_core_keymem_U2023 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[972]), .Y(aes_core_keymem_n1461) );
  OAI2BB2X1 aes_core_keymem_U2022 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1100]), .Y(aes_core_keymem_n1462) );
  OAI2BB2X1 aes_core_keymem_U2021 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1228]), .Y(aes_core_keymem_n1463) );
  OAI2BB2X1 aes_core_keymem_U2020 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1356]), .Y(aes_core_keymem_n1464) );
  OAI2BB2X1 aes_core_keymem_U2019 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[971]), .Y(aes_core_keymem_n1473) );
  OAI2BB2X1 aes_core_keymem_U2018 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1099]), .Y(aes_core_keymem_n1474) );
  OAI2BB2X1 aes_core_keymem_U2017 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1227]), .Y(aes_core_keymem_n1475) );
  OAI2BB2X1 aes_core_keymem_U2016 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1355]), .Y(aes_core_keymem_n1476) );
  OAI2BB2X1 aes_core_keymem_U2015 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[970]), .Y(aes_core_keymem_n1485) );
  OAI2BB2X1 aes_core_keymem_U2014 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1098]), .Y(aes_core_keymem_n1486) );
  OAI2BB2X1 aes_core_keymem_U2013 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1226]), .Y(aes_core_keymem_n1487) );
  OAI2BB2X1 aes_core_keymem_U2012 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1354]), .Y(aes_core_keymem_n1488) );
  OAI2BB2X1 aes_core_keymem_U2011 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[969]), .Y(aes_core_keymem_n1497) );
  OAI2BB2X1 aes_core_keymem_U2010 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1097]), .Y(aes_core_keymem_n1498) );
  OAI2BB2X1 aes_core_keymem_U2009 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1225]), .Y(aes_core_keymem_n1499) );
  OAI2BB2X1 aes_core_keymem_U2008 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1353]), .Y(aes_core_keymem_n1500) );
  OAI2BB2X1 aes_core_keymem_U2007 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[968]), .Y(aes_core_keymem_n1509) );
  OAI2BB2X1 aes_core_keymem_U2006 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1096]), .Y(aes_core_keymem_n1510) );
  OAI2BB2X1 aes_core_keymem_U2005 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1224]), .Y(aes_core_keymem_n1511) );
  OAI2BB2X1 aes_core_keymem_U2004 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1352]), .Y(aes_core_keymem_n1512) );
  OAI2BB2X1 aes_core_keymem_U2003 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[967]), .Y(aes_core_keymem_n1521) );
  OAI2BB2X1 aes_core_keymem_U2002 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1095]), .Y(aes_core_keymem_n1522) );
  OAI2BB2X1 aes_core_keymem_U2001 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1223]), .Y(aes_core_keymem_n1523) );
  OAI2BB2X1 aes_core_keymem_U2000 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1351]), .Y(aes_core_keymem_n1524) );
  OAI2BB2X1 aes_core_keymem_U1999 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[966]), .Y(aes_core_keymem_n1533) );
  OAI2BB2X1 aes_core_keymem_U1998 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1094]), .Y(aes_core_keymem_n1534) );
  OAI2BB2X1 aes_core_keymem_U1997 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1222]), .Y(aes_core_keymem_n1535) );
  OAI2BB2X1 aes_core_keymem_U1996 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1350]), .Y(aes_core_keymem_n1536) );
  OAI2BB2X1 aes_core_keymem_U1995 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[965]), .Y(aes_core_keymem_n1545) );
  OAI2BB2X1 aes_core_keymem_U1994 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1093]), .Y(aes_core_keymem_n1546) );
  OAI2BB2X1 aes_core_keymem_U1993 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1221]), .Y(aes_core_keymem_n1547) );
  OAI2BB2X1 aes_core_keymem_U1992 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1349]), .Y(aes_core_keymem_n1548) );
  OAI2BB2X1 aes_core_keymem_U1991 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[964]), .Y(aes_core_keymem_n1557) );
  OAI2BB2X1 aes_core_keymem_U1990 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1092]), .Y(aes_core_keymem_n1558) );
  OAI2BB2X1 aes_core_keymem_U1989 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1220]), .Y(aes_core_keymem_n1559) );
  OAI2BB2X1 aes_core_keymem_U1988 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1348]), .Y(aes_core_keymem_n1560) );
  OAI2BB2X1 aes_core_keymem_U1987 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n2630), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[963]), .Y(aes_core_keymem_n1569) );
  OAI2BB2X1 aes_core_keymem_U1986 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n2614), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1091]), .Y(aes_core_keymem_n1570) );
  OAI2BB2X1 aes_core_keymem_U1985 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n2597), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1219]), .Y(aes_core_keymem_n1571) );
  OAI2BB2X1 aes_core_keymem_U1984 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n2510), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1347]), .Y(aes_core_keymem_n1572) );
  OAI2BB2X1 aes_core_keymem_U1983 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[962]), .Y(aes_core_keymem_n1581) );
  OAI2BB2X1 aes_core_keymem_U1982 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1090]), .Y(aes_core_keymem_n1582) );
  OAI2BB2X1 aes_core_keymem_U1981 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1218]), .Y(aes_core_keymem_n1583) );
  OAI2BB2X1 aes_core_keymem_U1980 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1346]), .Y(aes_core_keymem_n1584) );
  OAI2BB2X1 aes_core_keymem_U1979 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[961]), .Y(aes_core_keymem_n1593) );
  OAI2BB2X1 aes_core_keymem_U1978 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1089]), .Y(aes_core_keymem_n1594) );
  OAI2BB2X1 aes_core_keymem_U1977 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1217]), .Y(aes_core_keymem_n1595) );
  OAI2BB2X1 aes_core_keymem_U1976 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1345]), .Y(aes_core_keymem_n1596) );
  OAI2BB2X1 aes_core_keymem_U1975 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[960]), .Y(aes_core_keymem_n1605) );
  OAI2BB2X1 aes_core_keymem_U1974 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1088]), .Y(aes_core_keymem_n1606) );
  OAI2BB2X1 aes_core_keymem_U1973 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1216]), .Y(aes_core_keymem_n1607) );
  OAI2BB2X1 aes_core_keymem_U1972 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1344]), .Y(aes_core_keymem_n1608) );
  OAI2BB2X1 aes_core_keymem_U1971 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[954]), .Y(aes_core_keymem_n1677) );
  OAI2BB2X1 aes_core_keymem_U1970 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1082]), .Y(aes_core_keymem_n1678) );
  OAI2BB2X1 aes_core_keymem_U1969 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1210]), .Y(aes_core_keymem_n1679) );
  OAI2BB2X1 aes_core_keymem_U1968 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1338]), .Y(aes_core_keymem_n1680) );
  OAI2BB2X1 aes_core_keymem_U1967 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[953]), .Y(aes_core_keymem_n1689) );
  OAI2BB2X1 aes_core_keymem_U1966 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1081]), .Y(aes_core_keymem_n1690) );
  OAI2BB2X1 aes_core_keymem_U1965 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1209]), .Y(aes_core_keymem_n1691) );
  OAI2BB2X1 aes_core_keymem_U1964 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1337]), .Y(aes_core_keymem_n1692) );
  OAI2BB2X1 aes_core_keymem_U1963 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[950]), .Y(aes_core_keymem_n1725) );
  OAI2BB2X1 aes_core_keymem_U1962 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1078]), .Y(aes_core_keymem_n1726) );
  OAI2BB2X1 aes_core_keymem_U1961 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1206]), .Y(aes_core_keymem_n1727) );
  OAI2BB2X1 aes_core_keymem_U1960 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1334]), .Y(aes_core_keymem_n1728) );
  OAI2BB2X1 aes_core_keymem_U1959 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[948]), .Y(aes_core_keymem_n1749) );
  OAI2BB2X1 aes_core_keymem_U1958 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1076]), .Y(aes_core_keymem_n1750) );
  OAI2BB2X1 aes_core_keymem_U1957 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1204]), .Y(aes_core_keymem_n1751) );
  OAI2BB2X1 aes_core_keymem_U1956 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1332]), .Y(aes_core_keymem_n1752) );
  OAI2BB2X1 aes_core_keymem_U1955 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[947]), .Y(aes_core_keymem_n1761) );
  OAI2BB2X1 aes_core_keymem_U1954 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1075]), .Y(aes_core_keymem_n1762) );
  OAI2BB2X1 aes_core_keymem_U1953 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1203]), .Y(aes_core_keymem_n1763) );
  OAI2BB2X1 aes_core_keymem_U1952 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1331]), .Y(aes_core_keymem_n1764) );
  OAI2BB2X1 aes_core_keymem_U1951 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[946]), .Y(aes_core_keymem_n1773) );
  OAI2BB2X1 aes_core_keymem_U1950 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1074]), .Y(aes_core_keymem_n1774) );
  OAI2BB2X1 aes_core_keymem_U1949 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1202]), .Y(aes_core_keymem_n1775) );
  OAI2BB2X1 aes_core_keymem_U1948 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1330]), .Y(aes_core_keymem_n1776) );
  OAI2BB2X1 aes_core_keymem_U1947 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[945]), .Y(aes_core_keymem_n1785) );
  OAI2BB2X1 aes_core_keymem_U1946 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1073]), .Y(aes_core_keymem_n1786) );
  OAI2BB2X1 aes_core_keymem_U1945 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1201]), .Y(aes_core_keymem_n1787) );
  OAI2BB2X1 aes_core_keymem_U1944 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1329]), .Y(aes_core_keymem_n1788) );
  OAI2BB2X1 aes_core_keymem_U1943 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[944]), .Y(aes_core_keymem_n1797) );
  OAI2BB2X1 aes_core_keymem_U1942 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1072]), .Y(aes_core_keymem_n1798) );
  OAI2BB2X1 aes_core_keymem_U1941 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1200]), .Y(aes_core_keymem_n1799) );
  OAI2BB2X1 aes_core_keymem_U1940 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1328]), .Y(aes_core_keymem_n1800) );
  OAI2BB2X1 aes_core_keymem_U1939 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2634), .A1N(
        aes_core_keymem_key_mem[938]), .Y(aes_core_keymem_n1869) );
  OAI2BB2X1 aes_core_keymem_U1938 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1066]), .Y(aes_core_keymem_n1870) );
  OAI2BB2X1 aes_core_keymem_U1937 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1194]), .Y(aes_core_keymem_n1871) );
  OAI2BB2X1 aes_core_keymem_U1936 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1322]), .Y(aes_core_keymem_n1872) );
  OAI2BB2X1 aes_core_keymem_U1935 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[937]), .Y(aes_core_keymem_n1881) );
  OAI2BB2X1 aes_core_keymem_U1934 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1065]), .Y(aes_core_keymem_n1882) );
  OAI2BB2X1 aes_core_keymem_U1933 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1193]), .Y(aes_core_keymem_n1883) );
  OAI2BB2X1 aes_core_keymem_U1932 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1321]), .Y(aes_core_keymem_n1884) );
  OAI2BB2X1 aes_core_keymem_U1931 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[934]), .Y(aes_core_keymem_n1917) );
  OAI2BB2X1 aes_core_keymem_U1930 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1062]), .Y(aes_core_keymem_n1918) );
  OAI2BB2X1 aes_core_keymem_U1929 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1190]), .Y(aes_core_keymem_n1919) );
  OAI2BB2X1 aes_core_keymem_U1928 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1318]), .Y(aes_core_keymem_n1920) );
  OAI2BB2X1 aes_core_keymem_U1927 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[933]), .Y(aes_core_keymem_n1929) );
  OAI2BB2X1 aes_core_keymem_U1926 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1061]), .Y(aes_core_keymem_n1930) );
  OAI2BB2X1 aes_core_keymem_U1925 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1189]), .Y(aes_core_keymem_n1931) );
  OAI2BB2X1 aes_core_keymem_U1924 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1317]), .Y(aes_core_keymem_n1932) );
  OAI2BB2X1 aes_core_keymem_U1923 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[932]), .Y(aes_core_keymem_n1941) );
  OAI2BB2X1 aes_core_keymem_U1922 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1060]), .Y(aes_core_keymem_n1942) );
  OAI2BB2X1 aes_core_keymem_U1921 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1188]), .Y(aes_core_keymem_n1943) );
  OAI2BB2X1 aes_core_keymem_U1920 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1316]), .Y(aes_core_keymem_n1944) );
  OAI2BB2X1 aes_core_keymem_U1919 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[931]), .Y(aes_core_keymem_n1953) );
  OAI2BB2X1 aes_core_keymem_U1918 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1059]), .Y(aes_core_keymem_n1954) );
  OAI2BB2X1 aes_core_keymem_U1917 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1187]), .Y(aes_core_keymem_n1955) );
  OAI2BB2X1 aes_core_keymem_U1916 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1315]), .Y(aes_core_keymem_n1956) );
  OAI2BB2X1 aes_core_keymem_U1915 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[930]), .Y(aes_core_keymem_n1965) );
  OAI2BB2X1 aes_core_keymem_U1914 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1058]), .Y(aes_core_keymem_n1966) );
  OAI2BB2X1 aes_core_keymem_U1913 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1186]), .Y(aes_core_keymem_n1967) );
  OAI2BB2X1 aes_core_keymem_U1912 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1314]), .Y(aes_core_keymem_n1968) );
  OAI2BB2X1 aes_core_keymem_U1911 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[929]), .Y(aes_core_keymem_n1977) );
  OAI2BB2X1 aes_core_keymem_U1910 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1057]), .Y(aes_core_keymem_n1978) );
  OAI2BB2X1 aes_core_keymem_U1909 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1185]), .Y(aes_core_keymem_n1979) );
  OAI2BB2X1 aes_core_keymem_U1908 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1313]), .Y(aes_core_keymem_n1980) );
  OAI2BB2X1 aes_core_keymem_U1907 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[928]), .Y(aes_core_keymem_n1989) );
  OAI2BB2X1 aes_core_keymem_U1906 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1056]), .Y(aes_core_keymem_n1990) );
  OAI2BB2X1 aes_core_keymem_U1905 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1184]), .Y(aes_core_keymem_n1991) );
  OAI2BB2X1 aes_core_keymem_U1904 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1312]), .Y(aes_core_keymem_n1992) );
  OAI2BB2X1 aes_core_keymem_U1903 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[912]), .Y(aes_core_keymem_n2181) );
  OAI2BB2X1 aes_core_keymem_U1902 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1040]), .Y(aes_core_keymem_n2182) );
  OAI2BB2X1 aes_core_keymem_U1901 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1168]), .Y(aes_core_keymem_n2183) );
  OAI2BB2X1 aes_core_keymem_U1900 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1296]), .Y(aes_core_keymem_n2184) );
  OAI2BB2X1 aes_core_keymem_U1899 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[901]), .Y(aes_core_keymem_n2313) );
  OAI2BB2X1 aes_core_keymem_U1898 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1029]), .Y(aes_core_keymem_n2314) );
  OAI2BB2X1 aes_core_keymem_U1897 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1157]), .Y(aes_core_keymem_n2315) );
  OAI2BB2X1 aes_core_keymem_U1896 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1285]), .Y(aes_core_keymem_n2316) );
  OAI2BB2X1 aes_core_keymem_U1895 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[897]), .Y(aes_core_keymem_n2361) );
  OAI2BB2X1 aes_core_keymem_U1894 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1025]), .Y(aes_core_keymem_n2362) );
  OAI2BB2X1 aes_core_keymem_U1893 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1153]), .Y(aes_core_keymem_n2363) );
  OAI2BB2X1 aes_core_keymem_U1892 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1281]), .Y(aes_core_keymem_n2364) );
  OAI2BB2X1 aes_core_keymem_U1891 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n2640), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[915]), .Y(aes_core_keymem_n2145) );
  OAI2BB2X1 aes_core_keymem_U1890 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n2623), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1043]), .Y(aes_core_keymem_n2146) );
  OAI2BB2X1 aes_core_keymem_U1889 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n2606), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1171]), .Y(aes_core_keymem_n2147) );
  OAI2BB2X1 aes_core_keymem_U1888 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1299]), .Y(aes_core_keymem_n2148) );
  OAI2BB2X1 aes_core_keymem_U1887 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n2638), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[914]), .Y(aes_core_keymem_n2157) );
  OAI2BB2X1 aes_core_keymem_U1886 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n2620), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1042]), .Y(aes_core_keymem_n2158) );
  OAI2BB2X1 aes_core_keymem_U1885 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n2603), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1170]), .Y(aes_core_keymem_n2159) );
  OAI2BB2X1 aes_core_keymem_U1884 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1298]), .Y(aes_core_keymem_n2160) );
  AOI22X1 aes_core_keymem_U1883 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n561), .B0(Din[254]), .B1(aes_core_keymem_n2522), .Y(
        aes_core_keymem_n560) );
  BUFX3 aes_core_keymem_U1882 ( .A(aes_core_keymem_n560), .Y(
        aes_core_keymem_n2504) );
  AOI22X1 aes_core_keymem_U1881 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n563), .B0(Din[253]), .B1(aes_core_keymem_n2523), .Y(
        aes_core_keymem_n562) );
  BUFX3 aes_core_keymem_U1880 ( .A(aes_core_keymem_n562), .Y(
        aes_core_keymem_n2503) );
  AOI22X1 aes_core_keymem_U1879 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n565), .B0(Din[252]), .B1(aes_core_keymem_n2523), .Y(
        aes_core_keymem_n564) );
  BUFX3 aes_core_keymem_U1878 ( .A(aes_core_keymem_n564), .Y(
        aes_core_keymem_n2502) );
  AOI22X1 aes_core_keymem_U1877 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n567), .B0(Din[251]), .B1(aes_core_keymem_n2524), .Y(
        aes_core_keymem_n566) );
  BUFX3 aes_core_keymem_U1876 ( .A(aes_core_keymem_n566), .Y(
        aes_core_keymem_n2501) );
  AOI22X1 aes_core_keymem_U1875 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n569), .B0(Din[250]), .B1(aes_core_keymem_n2524), .Y(
        aes_core_keymem_n568) );
  BUFX3 aes_core_keymem_U1874 ( .A(aes_core_keymem_n568), .Y(
        aes_core_keymem_n2500) );
  AOI22X1 aes_core_keymem_U1873 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n571), .B0(Din[249]), .B1(aes_core_keymem_n2525), .Y(
        aes_core_keymem_n570) );
  BUFX3 aes_core_keymem_U1872 ( .A(aes_core_keymem_n570), .Y(
        aes_core_keymem_n2499) );
  AOI22X1 aes_core_keymem_U1871 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n573), .B0(Din[248]), .B1(aes_core_keymem_n2525), .Y(
        aes_core_keymem_n572) );
  BUFX3 aes_core_keymem_U1870 ( .A(aes_core_keymem_n572), .Y(
        aes_core_keymem_n2498) );
  AOI22X1 aes_core_keymem_U1869 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n575), .B0(Din[247]), .B1(aes_core_keymem_n2526), .Y(
        aes_core_keymem_n574) );
  BUFX3 aes_core_keymem_U1868 ( .A(aes_core_keymem_n574), .Y(
        aes_core_keymem_n2497) );
  AOI22X1 aes_core_keymem_U1867 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n577), .B0(Din[246]), .B1(aes_core_keymem_n2526), .Y(
        aes_core_keymem_n576) );
  BUFX3 aes_core_keymem_U1866 ( .A(aes_core_keymem_n576), .Y(
        aes_core_keymem_n2496) );
  AOI22X1 aes_core_keymem_U1865 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n579), .B0(Din[245]), .B1(aes_core_keymem_n2527), .Y(
        aes_core_keymem_n578) );
  BUFX3 aes_core_keymem_U1864 ( .A(aes_core_keymem_n578), .Y(
        aes_core_keymem_n2495) );
  AOI22X1 aes_core_keymem_U1863 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n581), .B0(Din[244]), .B1(aes_core_keymem_n2527), .Y(
        aes_core_keymem_n580) );
  BUFX3 aes_core_keymem_U1862 ( .A(aes_core_keymem_n580), .Y(
        aes_core_keymem_n2494) );
  AOI22X1 aes_core_keymem_U1861 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n583), .B0(Din[243]), .B1(aes_core_keymem_n2528), .Y(
        aes_core_keymem_n582) );
  BUFX3 aes_core_keymem_U1860 ( .A(aes_core_keymem_n582), .Y(
        aes_core_keymem_n2493) );
  AOI22X1 aes_core_keymem_U1859 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n585), .B0(Din[242]), .B1(aes_core_keymem_n2528), .Y(
        aes_core_keymem_n584) );
  BUFX3 aes_core_keymem_U1858 ( .A(aes_core_keymem_n584), .Y(
        aes_core_keymem_n2492) );
  AOI22X1 aes_core_keymem_U1857 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n587), .B0(Din[241]), .B1(aes_core_keymem_n2529), .Y(
        aes_core_keymem_n586) );
  BUFX3 aes_core_keymem_U1856 ( .A(aes_core_keymem_n586), .Y(
        aes_core_keymem_n2491) );
  AOI22X1 aes_core_keymem_U1855 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n589), .B0(Din[240]), .B1(aes_core_keymem_n2529), .Y(
        aes_core_keymem_n588) );
  BUFX3 aes_core_keymem_U1854 ( .A(aes_core_keymem_n588), .Y(
        aes_core_keymem_n2490) );
  AOI22X1 aes_core_keymem_U1853 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n593), .B0(Din[238]), .B1(aes_core_keymem_n2530), .Y(
        aes_core_keymem_n592) );
  BUFX3 aes_core_keymem_U1852 ( .A(aes_core_keymem_n592), .Y(
        aes_core_keymem_n2488) );
  AOI22X1 aes_core_keymem_U1851 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n595), .B0(Din[237]), .B1(aes_core_keymem_n2531), .Y(
        aes_core_keymem_n594) );
  BUFX3 aes_core_keymem_U1850 ( .A(aes_core_keymem_n594), .Y(
        aes_core_keymem_n2487) );
  AOI22X1 aes_core_keymem_U1849 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n597), .B0(Din[236]), .B1(aes_core_keymem_n2531), .Y(
        aes_core_keymem_n596) );
  BUFX3 aes_core_keymem_U1848 ( .A(aes_core_keymem_n596), .Y(
        aes_core_keymem_n2486) );
  AOI22X1 aes_core_keymem_U1847 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n599), .B0(Din[235]), .B1(aes_core_keymem_n2525), .Y(
        aes_core_keymem_n598) );
  BUFX3 aes_core_keymem_U1846 ( .A(aes_core_keymem_n598), .Y(
        aes_core_keymem_n2485) );
  AOI22X1 aes_core_keymem_U1845 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n601), .B0(Din[234]), .B1(aes_core_keymem_n2526), .Y(
        aes_core_keymem_n600) );
  BUFX3 aes_core_keymem_U1844 ( .A(aes_core_keymem_n600), .Y(
        aes_core_keymem_n2484) );
  AOI22X1 aes_core_keymem_U1843 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n603), .B0(Din[233]), .B1(aes_core_keymem_n2532), .Y(
        aes_core_keymem_n602) );
  BUFX3 aes_core_keymem_U1842 ( .A(aes_core_keymem_n602), .Y(
        aes_core_keymem_n2483) );
  AOI22X1 aes_core_keymem_U1841 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n605), .B0(Din[232]), .B1(aes_core_keymem_n2532), .Y(
        aes_core_keymem_n604) );
  BUFX3 aes_core_keymem_U1840 ( .A(aes_core_keymem_n604), .Y(
        aes_core_keymem_n2482) );
  AOI22X1 aes_core_keymem_U1839 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n607), .B0(Din[231]), .B1(aes_core_keymem_n2533), .Y(
        aes_core_keymem_n606) );
  BUFX3 aes_core_keymem_U1838 ( .A(aes_core_keymem_n606), .Y(
        aes_core_keymem_n2481) );
  AOI22X1 aes_core_keymem_U1837 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n609), .B0(Din[230]), .B1(aes_core_keymem_n2533), .Y(
        aes_core_keymem_n608) );
  BUFX3 aes_core_keymem_U1836 ( .A(aes_core_keymem_n608), .Y(
        aes_core_keymem_n2480) );
  AOI22X1 aes_core_keymem_U1835 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n611), .B0(Din[229]), .B1(aes_core_keymem_n2534), .Y(
        aes_core_keymem_n610) );
  BUFX3 aes_core_keymem_U1834 ( .A(aes_core_keymem_n610), .Y(
        aes_core_keymem_n2479) );
  AOI22X1 aes_core_keymem_U1833 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n613), .B0(Din[228]), .B1(aes_core_keymem_n2534), .Y(
        aes_core_keymem_n612) );
  BUFX3 aes_core_keymem_U1832 ( .A(aes_core_keymem_n612), .Y(
        aes_core_keymem_n2478) );
  AOI22X1 aes_core_keymem_U1831 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n615), .B0(Din[227]), .B1(aes_core_keymem_n2535), .Y(
        aes_core_keymem_n614) );
  BUFX3 aes_core_keymem_U1830 ( .A(aes_core_keymem_n614), .Y(
        aes_core_keymem_n2477) );
  AOI22X1 aes_core_keymem_U1829 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n617), .B0(Din[226]), .B1(aes_core_keymem_n2535), .Y(
        aes_core_keymem_n616) );
  BUFX3 aes_core_keymem_U1828 ( .A(aes_core_keymem_n616), .Y(
        aes_core_keymem_n2476) );
  AOI22X1 aes_core_keymem_U1827 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n619), .B0(Din[225]), .B1(aes_core_keymem_n2536), .Y(
        aes_core_keymem_n618) );
  BUFX3 aes_core_keymem_U1826 ( .A(aes_core_keymem_n618), .Y(
        aes_core_keymem_n2475) );
  AOI22X1 aes_core_keymem_U1825 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n621), .B0(Din[224]), .B1(aes_core_keymem_n2536), .Y(
        aes_core_keymem_n620) );
  BUFX3 aes_core_keymem_U1824 ( .A(aes_core_keymem_n620), .Y(
        aes_core_keymem_n2474) );
  AOI22X1 aes_core_keymem_U1823 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n633), .B0(Din[218]), .B1(aes_core_keymem_n2541), .Y(
        aes_core_keymem_n632) );
  BUFX3 aes_core_keymem_U1822 ( .A(aes_core_keymem_n632), .Y(
        aes_core_keymem_n2468) );
  AOI22X1 aes_core_keymem_U1821 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n635), .B0(Din[217]), .B1(aes_core_keymem_n2539), .Y(
        aes_core_keymem_n634) );
  BUFX3 aes_core_keymem_U1820 ( .A(aes_core_keymem_n634), .Y(
        aes_core_keymem_n2467) );
  AOI22X1 aes_core_keymem_U1819 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n641), .B0(Din[214]), .B1(aes_core_keymem_n2540), .Y(
        aes_core_keymem_n640) );
  BUFX3 aes_core_keymem_U1818 ( .A(aes_core_keymem_n640), .Y(
        aes_core_keymem_n2464) );
  AOI22X1 aes_core_keymem_U1817 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n645), .B0(Din[212]), .B1(aes_core_keymem_n2541), .Y(
        aes_core_keymem_n644) );
  BUFX3 aes_core_keymem_U1816 ( .A(aes_core_keymem_n644), .Y(
        aes_core_keymem_n2462) );
  AOI22X1 aes_core_keymem_U1815 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n647), .B0(Din[211]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n646) );
  BUFX3 aes_core_keymem_U1814 ( .A(aes_core_keymem_n646), .Y(
        aes_core_keymem_n2461) );
  AOI22X1 aes_core_keymem_U1813 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n649), .B0(Din[210]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n648) );
  BUFX3 aes_core_keymem_U1812 ( .A(aes_core_keymem_n648), .Y(
        aes_core_keymem_n2460) );
  AOI22X1 aes_core_keymem_U1811 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n651), .B0(Din[209]), .B1(aes_core_keymem_n2542), .Y(
        aes_core_keymem_n650) );
  BUFX3 aes_core_keymem_U1810 ( .A(aes_core_keymem_n650), .Y(
        aes_core_keymem_n2459) );
  AOI22X1 aes_core_keymem_U1809 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n653), .B0(Din[208]), .B1(aes_core_keymem_n2542), .Y(
        aes_core_keymem_n652) );
  BUFX3 aes_core_keymem_U1808 ( .A(aes_core_keymem_n652), .Y(
        aes_core_keymem_n2458) );
  AOI22X1 aes_core_keymem_U1807 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n657), .B0(Din[206]), .B1(aes_core_keymem_n2543), .Y(
        aes_core_keymem_n656) );
  BUFX3 aes_core_keymem_U1806 ( .A(aes_core_keymem_n656), .Y(
        aes_core_keymem_n2456) );
  AOI22X1 aes_core_keymem_U1805 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n665), .B0(Din[202]), .B1(aes_core_keymem_n2545), .Y(
        aes_core_keymem_n664) );
  BUFX3 aes_core_keymem_U1804 ( .A(aes_core_keymem_n664), .Y(
        aes_core_keymem_n2452) );
  AOI22X1 aes_core_keymem_U1803 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n667), .B0(Din[201]), .B1(aes_core_keymem_n2546), .Y(
        aes_core_keymem_n666) );
  BUFX3 aes_core_keymem_U1802 ( .A(aes_core_keymem_n666), .Y(
        aes_core_keymem_n2451) );
  AOI22X1 aes_core_keymem_U1801 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n673), .B0(Din[198]), .B1(aes_core_keymem_n2547), .Y(
        aes_core_keymem_n672) );
  BUFX3 aes_core_keymem_U1800 ( .A(aes_core_keymem_n672), .Y(
        aes_core_keymem_n2448) );
  AOI22X1 aes_core_keymem_U1799 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n675), .B0(Din[197]), .B1(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n674) );
  BUFX3 aes_core_keymem_U1798 ( .A(aes_core_keymem_n674), .Y(
        aes_core_keymem_n2447) );
  AOI22X1 aes_core_keymem_U1797 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n677), .B0(Din[196]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n676) );
  BUFX3 aes_core_keymem_U1796 ( .A(aes_core_keymem_n676), .Y(
        aes_core_keymem_n2446) );
  AOI22X1 aes_core_keymem_U1795 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n679), .B0(Din[195]), .B1(aes_core_keymem_n2548), .Y(
        aes_core_keymem_n678) );
  BUFX3 aes_core_keymem_U1794 ( .A(aes_core_keymem_n678), .Y(
        aes_core_keymem_n2445) );
  AOI22X1 aes_core_keymem_U1793 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n681), .B0(Din[194]), .B1(aes_core_keymem_n2548), .Y(
        aes_core_keymem_n680) );
  BUFX3 aes_core_keymem_U1792 ( .A(aes_core_keymem_n680), .Y(
        aes_core_keymem_n2444) );
  AOI22X1 aes_core_keymem_U1791 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n683), .B0(Din[193]), .B1(aes_core_keymem_n2549), .Y(
        aes_core_keymem_n682) );
  BUFX3 aes_core_keymem_U1790 ( .A(aes_core_keymem_n682), .Y(
        aes_core_keymem_n2443) );
  AOI22X1 aes_core_keymem_U1789 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n685), .B0(Din[192]), .B1(aes_core_keymem_n2549), .Y(
        aes_core_keymem_n684) );
  BUFX3 aes_core_keymem_U1788 ( .A(aes_core_keymem_n684), .Y(
        aes_core_keymem_n2442) );
  AOI22X1 aes_core_keymem_U1787 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n711), .B0(Din[179]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n710) );
  BUFX3 aes_core_keymem_U1786 ( .A(aes_core_keymem_n710), .Y(
        aes_core_keymem_n2429) );
  AOI22X1 aes_core_keymem_U1785 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n713), .B0(Din[178]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n712) );
  BUFX3 aes_core_keymem_U1784 ( .A(aes_core_keymem_n712), .Y(
        aes_core_keymem_n2428) );
  AOI22X1 aes_core_keymem_U1783 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n747), .B0(Din[161]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n746) );
  BUFX3 aes_core_keymem_U1782 ( .A(aes_core_keymem_n746), .Y(
        aes_core_keymem_n2411) );
  OAI2BB2X1 aes_core_keymem_U1781 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n2628), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[991]), .Y(aes_core_keymem_n1233) );
  OAI2BB2X1 aes_core_keymem_U1780 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n2612), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1119]), .Y(aes_core_keymem_n1234) );
  OAI2BB2X1 aes_core_keymem_U1779 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n2595), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1247]), .Y(aes_core_keymem_n1235) );
  OAI2BB2X1 aes_core_keymem_U1778 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n2508), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1375]), .Y(aes_core_keymem_n1236) );
  OAI2BB2X1 aes_core_keymem_U1777 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n2629), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[975]), .Y(aes_core_keymem_n1425) );
  OAI2BB2X1 aes_core_keymem_U1776 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n2613), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1103]), .Y(aes_core_keymem_n1426) );
  OAI2BB2X1 aes_core_keymem_U1775 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n2596), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1231]), .Y(aes_core_keymem_n1427) );
  OAI2BB2X1 aes_core_keymem_U1774 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n2509), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1359]), .Y(aes_core_keymem_n1428) );
  OAI2BB2X1 aes_core_keymem_U1773 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[959]), .Y(aes_core_keymem_n1617) );
  OAI2BB2X1 aes_core_keymem_U1772 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1087]), .Y(aes_core_keymem_n1618) );
  OAI2BB2X1 aes_core_keymem_U1771 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1215]), .Y(aes_core_keymem_n1619) );
  OAI2BB2X1 aes_core_keymem_U1770 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1343]), .Y(aes_core_keymem_n1620) );
  OAI2BB2X1 aes_core_keymem_U1769 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[958]), .Y(aes_core_keymem_n1629) );
  OAI2BB2X1 aes_core_keymem_U1768 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1086]), .Y(aes_core_keymem_n1630) );
  OAI2BB2X1 aes_core_keymem_U1767 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1214]), .Y(aes_core_keymem_n1631) );
  OAI2BB2X1 aes_core_keymem_U1766 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1342]), .Y(aes_core_keymem_n1632) );
  OAI2BB2X1 aes_core_keymem_U1765 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[957]), .Y(aes_core_keymem_n1641) );
  OAI2BB2X1 aes_core_keymem_U1764 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1085]), .Y(aes_core_keymem_n1642) );
  OAI2BB2X1 aes_core_keymem_U1763 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1213]), .Y(aes_core_keymem_n1643) );
  OAI2BB2X1 aes_core_keymem_U1762 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1341]), .Y(aes_core_keymem_n1644) );
  OAI2BB2X1 aes_core_keymem_U1761 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[956]), .Y(aes_core_keymem_n1653) );
  OAI2BB2X1 aes_core_keymem_U1760 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1084]), .Y(aes_core_keymem_n1654) );
  OAI2BB2X1 aes_core_keymem_U1759 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1212]), .Y(aes_core_keymem_n1655) );
  OAI2BB2X1 aes_core_keymem_U1758 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1340]), .Y(aes_core_keymem_n1656) );
  OAI2BB2X1 aes_core_keymem_U1757 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[955]), .Y(aes_core_keymem_n1665) );
  OAI2BB2X1 aes_core_keymem_U1756 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1083]), .Y(aes_core_keymem_n1666) );
  OAI2BB2X1 aes_core_keymem_U1755 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1211]), .Y(aes_core_keymem_n1667) );
  OAI2BB2X1 aes_core_keymem_U1754 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1339]), .Y(aes_core_keymem_n1668) );
  OAI2BB2X1 aes_core_keymem_U1753 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[952]), .Y(aes_core_keymem_n1701) );
  OAI2BB2X1 aes_core_keymem_U1752 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1080]), .Y(aes_core_keymem_n1702) );
  OAI2BB2X1 aes_core_keymem_U1751 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1208]), .Y(aes_core_keymem_n1703) );
  OAI2BB2X1 aes_core_keymem_U1750 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1336]), .Y(aes_core_keymem_n1704) );
  OAI2BB2X1 aes_core_keymem_U1749 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n2631), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[951]), .Y(aes_core_keymem_n1713) );
  OAI2BB2X1 aes_core_keymem_U1748 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n2615), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1079]), .Y(aes_core_keymem_n1714) );
  OAI2BB2X1 aes_core_keymem_U1747 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n2598), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1207]), .Y(aes_core_keymem_n1715) );
  OAI2BB2X1 aes_core_keymem_U1746 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n2511), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1335]), .Y(aes_core_keymem_n1716) );
  OAI2BB2X1 aes_core_keymem_U1745 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[949]), .Y(aes_core_keymem_n1737) );
  OAI2BB2X1 aes_core_keymem_U1744 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1077]), .Y(aes_core_keymem_n1738) );
  OAI2BB2X1 aes_core_keymem_U1743 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1205]), .Y(aes_core_keymem_n1739) );
  OAI2BB2X1 aes_core_keymem_U1742 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1333]), .Y(aes_core_keymem_n1740) );
  OAI2BB2X1 aes_core_keymem_U1741 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[943]), .Y(aes_core_keymem_n1809) );
  OAI2BB2X1 aes_core_keymem_U1740 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1071]), .Y(aes_core_keymem_n1810) );
  OAI2BB2X1 aes_core_keymem_U1739 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1199]), .Y(aes_core_keymem_n1811) );
  OAI2BB2X1 aes_core_keymem_U1738 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1327]), .Y(aes_core_keymem_n1812) );
  OAI2BB2X1 aes_core_keymem_U1737 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[942]), .Y(aes_core_keymem_n1821) );
  OAI2BB2X1 aes_core_keymem_U1736 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1070]), .Y(aes_core_keymem_n1822) );
  OAI2BB2X1 aes_core_keymem_U1735 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1198]), .Y(aes_core_keymem_n1823) );
  OAI2BB2X1 aes_core_keymem_U1734 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1326]), .Y(aes_core_keymem_n1824) );
  OAI2BB2X1 aes_core_keymem_U1733 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[941]), .Y(aes_core_keymem_n1833) );
  OAI2BB2X1 aes_core_keymem_U1732 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1069]), .Y(aes_core_keymem_n1834) );
  OAI2BB2X1 aes_core_keymem_U1731 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1197]), .Y(aes_core_keymem_n1835) );
  OAI2BB2X1 aes_core_keymem_U1730 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1325]), .Y(aes_core_keymem_n1836) );
  OAI2BB2X1 aes_core_keymem_U1729 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2632), .A1N(
        aes_core_keymem_key_mem[940]), .Y(aes_core_keymem_n1845) );
  OAI2BB2X1 aes_core_keymem_U1728 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1068]), .Y(aes_core_keymem_n1846) );
  OAI2BB2X1 aes_core_keymem_U1727 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1196]), .Y(aes_core_keymem_n1847) );
  OAI2BB2X1 aes_core_keymem_U1726 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1324]), .Y(aes_core_keymem_n1848) );
  OAI2BB2X1 aes_core_keymem_U1725 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[939]), .Y(aes_core_keymem_n1857) );
  OAI2BB2X1 aes_core_keymem_U1724 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n2616), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1067]), .Y(aes_core_keymem_n1858) );
  OAI2BB2X1 aes_core_keymem_U1723 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n2599), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1195]), .Y(aes_core_keymem_n1859) );
  OAI2BB2X1 aes_core_keymem_U1722 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n2512), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1323]), .Y(aes_core_keymem_n1860) );
  OAI2BB2X1 aes_core_keymem_U1721 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[936]), .Y(aes_core_keymem_n1893) );
  OAI2BB2X1 aes_core_keymem_U1720 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1064]), .Y(aes_core_keymem_n1894) );
  OAI2BB2X1 aes_core_keymem_U1719 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1192]), .Y(aes_core_keymem_n1895) );
  OAI2BB2X1 aes_core_keymem_U1718 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1320]), .Y(aes_core_keymem_n1896) );
  OAI2BB2X1 aes_core_keymem_U1717 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[935]), .Y(aes_core_keymem_n1905) );
  OAI2BB2X1 aes_core_keymem_U1716 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1063]), .Y(aes_core_keymem_n1906) );
  OAI2BB2X1 aes_core_keymem_U1715 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1191]), .Y(aes_core_keymem_n1907) );
  OAI2BB2X1 aes_core_keymem_U1714 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1319]), .Y(aes_core_keymem_n1908) );
  OAI2BB2X1 aes_core_keymem_U1713 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[927]), .Y(aes_core_keymem_n2001) );
  OAI2BB2X1 aes_core_keymem_U1712 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1055]), .Y(aes_core_keymem_n2002) );
  OAI2BB2X1 aes_core_keymem_U1711 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1183]), .Y(aes_core_keymem_n2003) );
  OAI2BB2X1 aes_core_keymem_U1710 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1311]), .Y(aes_core_keymem_n2004) );
  OAI2BB2X1 aes_core_keymem_U1709 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2640), .A1N(
        aes_core_keymem_key_mem[926]), .Y(aes_core_keymem_n2013) );
  OAI2BB2X1 aes_core_keymem_U1708 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2623), .A1N(
        aes_core_keymem_key_mem[1054]), .Y(aes_core_keymem_n2014) );
  OAI2BB2X1 aes_core_keymem_U1707 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2606), .A1N(
        aes_core_keymem_key_mem[1182]), .Y(aes_core_keymem_n2015) );
  OAI2BB2X1 aes_core_keymem_U1706 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1310]), .Y(aes_core_keymem_n2016) );
  OAI2BB2X1 aes_core_keymem_U1705 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[925]), .Y(aes_core_keymem_n2025) );
  OAI2BB2X1 aes_core_keymem_U1704 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1053]), .Y(aes_core_keymem_n2026) );
  OAI2BB2X1 aes_core_keymem_U1703 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1181]), .Y(aes_core_keymem_n2027) );
  OAI2BB2X1 aes_core_keymem_U1702 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1309]), .Y(aes_core_keymem_n2028) );
  OAI2BB2X1 aes_core_keymem_U1701 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[924]), .Y(aes_core_keymem_n2037) );
  OAI2BB2X1 aes_core_keymem_U1700 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1052]), .Y(aes_core_keymem_n2038) );
  OAI2BB2X1 aes_core_keymem_U1699 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1180]), .Y(aes_core_keymem_n2039) );
  OAI2BB2X1 aes_core_keymem_U1698 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1308]), .Y(aes_core_keymem_n2040) );
  OAI2BB2X1 aes_core_keymem_U1697 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[923]), .Y(aes_core_keymem_n2049) );
  OAI2BB2X1 aes_core_keymem_U1696 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1051]), .Y(aes_core_keymem_n2050) );
  OAI2BB2X1 aes_core_keymem_U1695 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1179]), .Y(aes_core_keymem_n2051) );
  OAI2BB2X1 aes_core_keymem_U1694 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1307]), .Y(aes_core_keymem_n2052) );
  OAI2BB2X1 aes_core_keymem_U1693 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[922]), .Y(aes_core_keymem_n2061) );
  OAI2BB2X1 aes_core_keymem_U1692 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1050]), .Y(aes_core_keymem_n2062) );
  OAI2BB2X1 aes_core_keymem_U1691 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1178]), .Y(aes_core_keymem_n2063) );
  OAI2BB2X1 aes_core_keymem_U1690 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2520), .A1N(
        aes_core_keymem_key_mem[1306]), .Y(aes_core_keymem_n2064) );
  OAI2BB2X1 aes_core_keymem_U1689 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2639), .A1N(
        aes_core_keymem_key_mem[921]), .Y(aes_core_keymem_n2073) );
  OAI2BB2X1 aes_core_keymem_U1688 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1049]), .Y(aes_core_keymem_n2074) );
  OAI2BB2X1 aes_core_keymem_U1687 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1177]), .Y(aes_core_keymem_n2075) );
  OAI2BB2X1 aes_core_keymem_U1686 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2521), .A1N(
        aes_core_keymem_key_mem[1305]), .Y(aes_core_keymem_n2076) );
  OAI2BB2X1 aes_core_keymem_U1685 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[920]), .Y(aes_core_keymem_n2085) );
  OAI2BB2X1 aes_core_keymem_U1684 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1048]), .Y(aes_core_keymem_n2086) );
  OAI2BB2X1 aes_core_keymem_U1683 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1176]), .Y(aes_core_keymem_n2087) );
  OAI2BB2X1 aes_core_keymem_U1682 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1304]), .Y(aes_core_keymem_n2088) );
  OAI2BB2X1 aes_core_keymem_U1681 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[916]), .Y(aes_core_keymem_n2133) );
  OAI2BB2X1 aes_core_keymem_U1680 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1044]), .Y(aes_core_keymem_n2134) );
  OAI2BB2X1 aes_core_keymem_U1679 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1172]), .Y(aes_core_keymem_n2135) );
  OAI2BB2X1 aes_core_keymem_U1678 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1300]), .Y(aes_core_keymem_n2136) );
  OAI2BB2X1 aes_core_keymem_U1677 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[909]), .Y(aes_core_keymem_n2217) );
  OAI2BB2X1 aes_core_keymem_U1676 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1037]), .Y(aes_core_keymem_n2218) );
  OAI2BB2X1 aes_core_keymem_U1675 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1165]), .Y(aes_core_keymem_n2219) );
  OAI2BB2X1 aes_core_keymem_U1674 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1293]), .Y(aes_core_keymem_n2220) );
  OAI2BB2X1 aes_core_keymem_U1673 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[908]), .Y(aes_core_keymem_n2229) );
  OAI2BB2X1 aes_core_keymem_U1672 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1036]), .Y(aes_core_keymem_n2230) );
  OAI2BB2X1 aes_core_keymem_U1671 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1164]), .Y(aes_core_keymem_n2231) );
  OAI2BB2X1 aes_core_keymem_U1670 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1292]), .Y(aes_core_keymem_n2232) );
  OAI2BB2X1 aes_core_keymem_U1669 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[907]), .Y(aes_core_keymem_n2241) );
  OAI2BB2X1 aes_core_keymem_U1668 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1035]), .Y(aes_core_keymem_n2242) );
  OAI2BB2X1 aes_core_keymem_U1667 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1163]), .Y(aes_core_keymem_n2243) );
  OAI2BB2X1 aes_core_keymem_U1666 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1291]), .Y(aes_core_keymem_n2244) );
  OAI2BB2X1 aes_core_keymem_U1665 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[906]), .Y(aes_core_keymem_n2253) );
  OAI2BB2X1 aes_core_keymem_U1664 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n555), .A1N(
        aes_core_keymem_key_mem[1034]), .Y(aes_core_keymem_n2254) );
  OAI2BB2X1 aes_core_keymem_U1663 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n556), .A1N(
        aes_core_keymem_key_mem[1162]), .Y(aes_core_keymem_n2255) );
  OAI2BB2X1 aes_core_keymem_U1662 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1290]), .Y(aes_core_keymem_n2256) );
  OAI2BB2X1 aes_core_keymem_U1661 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[905]), .Y(aes_core_keymem_n2265) );
  OAI2BB2X1 aes_core_keymem_U1660 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2624), .A1N(
        aes_core_keymem_key_mem[1033]), .Y(aes_core_keymem_n2266) );
  OAI2BB2X1 aes_core_keymem_U1659 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2607), .A1N(
        aes_core_keymem_key_mem[1161]), .Y(aes_core_keymem_n2267) );
  OAI2BB2X1 aes_core_keymem_U1658 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1289]), .Y(aes_core_keymem_n2268) );
  OAI2BB2X1 aes_core_keymem_U1657 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n2634), .A0N(aes_core_keymem_n2636), .A1N(
        aes_core_keymem_key_mem[904]), .Y(aes_core_keymem_n2277) );
  OAI2BB2X1 aes_core_keymem_U1656 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n2619), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1032]), .Y(aes_core_keymem_n2278) );
  OAI2BB2X1 aes_core_keymem_U1655 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n2602), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1160]), .Y(aes_core_keymem_n2279) );
  OAI2BB2X1 aes_core_keymem_U1654 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n2515), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1288]), .Y(aes_core_keymem_n2280) );
  OAI2BB2X1 aes_core_keymem_U1653 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[903]), .Y(aes_core_keymem_n2289) );
  OAI2BB2X1 aes_core_keymem_U1652 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1031]), .Y(aes_core_keymem_n2290) );
  OAI2BB2X1 aes_core_keymem_U1651 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1159]), .Y(aes_core_keymem_n2291) );
  OAI2BB2X1 aes_core_keymem_U1650 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1287]), .Y(aes_core_keymem_n2292) );
  OAI2BB2X1 aes_core_keymem_U1649 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[902]), .Y(aes_core_keymem_n2301) );
  OAI2BB2X1 aes_core_keymem_U1648 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1030]), .Y(aes_core_keymem_n2302) );
  OAI2BB2X1 aes_core_keymem_U1647 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1158]), .Y(aes_core_keymem_n2303) );
  OAI2BB2X1 aes_core_keymem_U1646 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1286]), .Y(aes_core_keymem_n2304) );
  OAI2BB2X1 aes_core_keymem_U1645 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[900]), .Y(aes_core_keymem_n2325) );
  OAI2BB2X1 aes_core_keymem_U1644 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1028]), .Y(aes_core_keymem_n2326) );
  OAI2BB2X1 aes_core_keymem_U1643 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1156]), .Y(aes_core_keymem_n2327) );
  OAI2BB2X1 aes_core_keymem_U1642 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1284]), .Y(aes_core_keymem_n2328) );
  OAI2BB2X1 aes_core_keymem_U1641 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n2633), .A0N(aes_core_keymem_n2635), .A1N(
        aes_core_keymem_key_mem[899]), .Y(aes_core_keymem_n2337) );
  OAI2BB2X1 aes_core_keymem_U1640 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n2618), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1027]), .Y(aes_core_keymem_n2338) );
  OAI2BB2X1 aes_core_keymem_U1639 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n2601), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1155]), .Y(aes_core_keymem_n2339) );
  OAI2BB2X1 aes_core_keymem_U1638 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n2514), .A0N(aes_core_keymem_n2517), .A1N(
        aes_core_keymem_key_mem[1283]), .Y(aes_core_keymem_n2340) );
  OAI2BB2X1 aes_core_keymem_U1637 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[898]), .Y(aes_core_keymem_n2349) );
  OAI2BB2X1 aes_core_keymem_U1636 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2620), .A1N(
        aes_core_keymem_key_mem[1026]), .Y(aes_core_keymem_n2350) );
  OAI2BB2X1 aes_core_keymem_U1635 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2603), .A1N(
        aes_core_keymem_key_mem[1154]), .Y(aes_core_keymem_n2351) );
  OAI2BB2X1 aes_core_keymem_U1634 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2516), .A1N(
        aes_core_keymem_key_mem[1282]), .Y(aes_core_keymem_n2352) );
  OAI2BB2X1 aes_core_keymem_U1633 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n2632), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[896]), .Y(aes_core_keymem_n2373) );
  OAI2BB2X1 aes_core_keymem_U1632 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n2617), .A0N(aes_core_keymem_n2622), .A1N(
        aes_core_keymem_key_mem[1024]), .Y(aes_core_keymem_n2374) );
  OAI2BB2X1 aes_core_keymem_U1631 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n2600), .A0N(aes_core_keymem_n2605), .A1N(
        aes_core_keymem_key_mem[1152]), .Y(aes_core_keymem_n2375) );
  OAI2BB2X1 aes_core_keymem_U1630 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n2513), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1280]), .Y(aes_core_keymem_n2376) );
  OAI2BB2X1 aes_core_keymem_U1629 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n2635), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[919]), .Y(aes_core_keymem_n2097) );
  OAI2BB2X1 aes_core_keymem_U1628 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n2609), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1047]), .Y(aes_core_keymem_n2098) );
  OAI2BB2X1 aes_core_keymem_U1627 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n2592), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1175]), .Y(aes_core_keymem_n2099) );
  OAI2BB2X1 aes_core_keymem_U1626 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1303]), .Y(aes_core_keymem_n2100) );
  OAI2BB2X1 aes_core_keymem_U1625 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n2636), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[918]), .Y(aes_core_keymem_n2109) );
  OAI2BB2X1 aes_core_keymem_U1624 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n2620), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1046]), .Y(aes_core_keymem_n2110) );
  OAI2BB2X1 aes_core_keymem_U1623 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n2603), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1174]), .Y(aes_core_keymem_n2111) );
  OAI2BB2X1 aes_core_keymem_U1622 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1302]), .Y(aes_core_keymem_n2112) );
  OAI2BB2X1 aes_core_keymem_U1621 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n2637), .A0N(aes_core_keymem_n2638), .A1N(
        aes_core_keymem_key_mem[917]), .Y(aes_core_keymem_n2121) );
  OAI2BB2X1 aes_core_keymem_U1620 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n2609), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1045]), .Y(aes_core_keymem_n2122) );
  OAI2BB2X1 aes_core_keymem_U1619 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n2592), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1173]), .Y(aes_core_keymem_n2123) );
  OAI2BB2X1 aes_core_keymem_U1618 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2519), .A1N(
        aes_core_keymem_key_mem[1301]), .Y(aes_core_keymem_n2124) );
  OAI2BB2X1 aes_core_keymem_U1617 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n2639), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[913]), .Y(aes_core_keymem_n2169) );
  OAI2BB2X1 aes_core_keymem_U1616 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n2620), .A0N(aes_core_keymem_n2609), .A1N(
        aes_core_keymem_key_mem[1041]), .Y(aes_core_keymem_n2170) );
  OAI2BB2X1 aes_core_keymem_U1615 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n2603), .A0N(aes_core_keymem_n2592), .A1N(
        aes_core_keymem_key_mem[1169]), .Y(aes_core_keymem_n2171) );
  OAI2BB2X1 aes_core_keymem_U1614 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1297]), .Y(aes_core_keymem_n2172) );
  OAI2BB2X1 aes_core_keymem_U1613 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n2640), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[911]), .Y(aes_core_keymem_n2193) );
  OAI2BB2X1 aes_core_keymem_U1612 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n2609), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1039]), .Y(aes_core_keymem_n2194) );
  OAI2BB2X1 aes_core_keymem_U1611 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n2592), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1167]), .Y(aes_core_keymem_n2195) );
  OAI2BB2X1 aes_core_keymem_U1610 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1295]), .Y(aes_core_keymem_n2196) );
  OAI2BB2X1 aes_core_keymem_U1609 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n2638), .A0N(aes_core_keymem_n2637), .A1N(
        aes_core_keymem_key_mem[910]), .Y(aes_core_keymem_n2205) );
  OAI2BB2X1 aes_core_keymem_U1608 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n2620), .A0N(aes_core_keymem_n2621), .A1N(
        aes_core_keymem_key_mem[1038]), .Y(aes_core_keymem_n2206) );
  OAI2BB2X1 aes_core_keymem_U1607 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n2603), .A0N(aes_core_keymem_n2604), .A1N(
        aes_core_keymem_key_mem[1166]), .Y(aes_core_keymem_n2207) );
  OAI2BB2X1 aes_core_keymem_U1606 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n2516), .A0N(aes_core_keymem_n2518), .A1N(
        aes_core_keymem_key_mem[1294]), .Y(aes_core_keymem_n2208) );
  AOI22X1 aes_core_keymem_U1605 ( .A0(aes_core_keymem_n2581), .A1(
        aes_core_keymem_n558), .B0(Din[255]), .B1(aes_core_keymem_n2522), .Y(
        aes_core_keymem_n546) );
  BUFX3 aes_core_keymem_U1604 ( .A(aes_core_keymem_n546), .Y(
        aes_core_keymem_n2505) );
  AOI22X1 aes_core_keymem_U1603 ( .A0(aes_core_keymem_n2582), .A1(
        aes_core_keymem_n591), .B0(Din[239]), .B1(aes_core_keymem_n2530), .Y(
        aes_core_keymem_n590) );
  BUFX3 aes_core_keymem_U1602 ( .A(aes_core_keymem_n590), .Y(
        aes_core_keymem_n2489) );
  AOI22X1 aes_core_keymem_U1601 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n623), .B0(Din[223]), .B1(aes_core_keymem_n2537), .Y(
        aes_core_keymem_n622) );
  BUFX3 aes_core_keymem_U1600 ( .A(aes_core_keymem_n622), .Y(
        aes_core_keymem_n2473) );
  AOI22X1 aes_core_keymem_U1599 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n625), .B0(Din[222]), .B1(aes_core_keymem_n2537), .Y(
        aes_core_keymem_n624) );
  BUFX3 aes_core_keymem_U1598 ( .A(aes_core_keymem_n624), .Y(
        aes_core_keymem_n2472) );
  AOI22X1 aes_core_keymem_U1597 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n627), .B0(Din[221]), .B1(aes_core_keymem_n2538), .Y(
        aes_core_keymem_n626) );
  BUFX3 aes_core_keymem_U1596 ( .A(aes_core_keymem_n626), .Y(
        aes_core_keymem_n2471) );
  AOI22X1 aes_core_keymem_U1595 ( .A0(aes_core_keymem_n2583), .A1(
        aes_core_keymem_n629), .B0(Din[220]), .B1(aes_core_keymem_n2538), .Y(
        aes_core_keymem_n628) );
  BUFX3 aes_core_keymem_U1594 ( .A(aes_core_keymem_n628), .Y(
        aes_core_keymem_n2470) );
  AOI22X1 aes_core_keymem_U1593 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n631), .B0(Din[219]), .B1(aes_core_keymem_n2538), .Y(
        aes_core_keymem_n630) );
  BUFX3 aes_core_keymem_U1592 ( .A(aes_core_keymem_n630), .Y(
        aes_core_keymem_n2469) );
  AOI22X1 aes_core_keymem_U1591 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n637), .B0(Din[216]), .B1(aes_core_keymem_n2539), .Y(
        aes_core_keymem_n636) );
  BUFX3 aes_core_keymem_U1590 ( .A(aes_core_keymem_n636), .Y(
        aes_core_keymem_n2466) );
  AOI22X1 aes_core_keymem_U1589 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n639), .B0(Din[215]), .B1(aes_core_keymem_n2540), .Y(
        aes_core_keymem_n638) );
  BUFX3 aes_core_keymem_U1588 ( .A(aes_core_keymem_n638), .Y(
        aes_core_keymem_n2465) );
  AOI22X1 aes_core_keymem_U1587 ( .A0(aes_core_keymem_n2584), .A1(
        aes_core_keymem_n643), .B0(Din[213]), .B1(aes_core_keymem_n2541), .Y(
        aes_core_keymem_n642) );
  BUFX3 aes_core_keymem_U1586 ( .A(aes_core_keymem_n642), .Y(
        aes_core_keymem_n2463) );
  AOI22X1 aes_core_keymem_U1585 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n655), .B0(Din[207]), .B1(aes_core_keymem_n2543), .Y(
        aes_core_keymem_n654) );
  BUFX3 aes_core_keymem_U1584 ( .A(aes_core_keymem_n654), .Y(
        aes_core_keymem_n2457) );
  AOI22X1 aes_core_keymem_U1583 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n659), .B0(Din[205]), .B1(aes_core_keymem_n2544), .Y(
        aes_core_keymem_n658) );
  BUFX3 aes_core_keymem_U1582 ( .A(aes_core_keymem_n658), .Y(
        aes_core_keymem_n2455) );
  AOI22X1 aes_core_keymem_U1581 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n661), .B0(Din[204]), .B1(aes_core_keymem_n2544), .Y(
        aes_core_keymem_n660) );
  BUFX3 aes_core_keymem_U1580 ( .A(aes_core_keymem_n660), .Y(
        aes_core_keymem_n2454) );
  AOI22X1 aes_core_keymem_U1579 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n663), .B0(Din[203]), .B1(aes_core_keymem_n2545), .Y(
        aes_core_keymem_n662) );
  BUFX3 aes_core_keymem_U1578 ( .A(aes_core_keymem_n662), .Y(
        aes_core_keymem_n2453) );
  AOI22X1 aes_core_keymem_U1577 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n669), .B0(Din[200]), .B1(aes_core_keymem_n2546), .Y(
        aes_core_keymem_n668) );
  BUFX3 aes_core_keymem_U1576 ( .A(aes_core_keymem_n668), .Y(
        aes_core_keymem_n2450) );
  AOI22X1 aes_core_keymem_U1575 ( .A0(aes_core_keymem_n2585), .A1(
        aes_core_keymem_n671), .B0(Din[199]), .B1(aes_core_keymem_n2547), .Y(
        aes_core_keymem_n670) );
  BUFX3 aes_core_keymem_U1574 ( .A(aes_core_keymem_n670), .Y(
        aes_core_keymem_n2449) );
  AOI22X1 aes_core_keymem_U1573 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n689), .B0(Din[190]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n688) );
  BUFX3 aes_core_keymem_U1572 ( .A(aes_core_keymem_n688), .Y(
        aes_core_keymem_n2440) );
  AOI22X1 aes_core_keymem_U1571 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n691), .B0(Din[189]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n690) );
  BUFX3 aes_core_keymem_U1570 ( .A(aes_core_keymem_n690), .Y(
        aes_core_keymem_n2439) );
  AOI22X1 aes_core_keymem_U1569 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n693), .B0(Din[188]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n692) );
  BUFX3 aes_core_keymem_U1568 ( .A(aes_core_keymem_n692), .Y(
        aes_core_keymem_n2438) );
  AOI22X1 aes_core_keymem_U1567 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n695), .B0(Din[187]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n694) );
  BUFX3 aes_core_keymem_U1566 ( .A(aes_core_keymem_n694), .Y(
        aes_core_keymem_n2437) );
  AOI22X1 aes_core_keymem_U1565 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n697), .B0(Din[186]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n696) );
  BUFX3 aes_core_keymem_U1564 ( .A(aes_core_keymem_n696), .Y(
        aes_core_keymem_n2436) );
  AOI22X1 aes_core_keymem_U1563 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n699), .B0(Din[185]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n698) );
  BUFX3 aes_core_keymem_U1562 ( .A(aes_core_keymem_n698), .Y(
        aes_core_keymem_n2435) );
  AOI22X1 aes_core_keymem_U1561 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n701), .B0(Din[184]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n700) );
  BUFX3 aes_core_keymem_U1560 ( .A(aes_core_keymem_n700), .Y(
        aes_core_keymem_n2434) );
  AOI22X1 aes_core_keymem_U1559 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n703), .B0(Din[183]), .B1(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n702) );
  BUFX3 aes_core_keymem_U1558 ( .A(aes_core_keymem_n702), .Y(
        aes_core_keymem_n2433) );
  AOI22X1 aes_core_keymem_U1557 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n705), .B0(Din[182]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n704) );
  BUFX3 aes_core_keymem_U1556 ( .A(aes_core_keymem_n704), .Y(
        aes_core_keymem_n2432) );
  AOI22X1 aes_core_keymem_U1555 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n707), .B0(Din[181]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n706) );
  BUFX3 aes_core_keymem_U1554 ( .A(aes_core_keymem_n706), .Y(
        aes_core_keymem_n2431) );
  AOI22X1 aes_core_keymem_U1553 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n709), .B0(Din[180]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n708) );
  BUFX3 aes_core_keymem_U1552 ( .A(aes_core_keymem_n708), .Y(
        aes_core_keymem_n2430) );
  AOI22X1 aes_core_keymem_U1551 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n715), .B0(Din[177]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n714) );
  BUFX3 aes_core_keymem_U1550 ( .A(aes_core_keymem_n714), .Y(
        aes_core_keymem_n2427) );
  AOI22X1 aes_core_keymem_U1549 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n717), .B0(Din[176]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n716) );
  BUFX3 aes_core_keymem_U1548 ( .A(aes_core_keymem_n716), .Y(
        aes_core_keymem_n2426) );
  AOI22X1 aes_core_keymem_U1547 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n719), .B0(Din[175]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n718) );
  BUFX3 aes_core_keymem_U1546 ( .A(aes_core_keymem_n718), .Y(
        aes_core_keymem_n2425) );
  AOI22X1 aes_core_keymem_U1545 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n721), .B0(Din[174]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n720) );
  BUFX3 aes_core_keymem_U1544 ( .A(aes_core_keymem_n720), .Y(
        aes_core_keymem_n2424) );
  AOI22X1 aes_core_keymem_U1543 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n723), .B0(Din[173]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n722) );
  BUFX3 aes_core_keymem_U1542 ( .A(aes_core_keymem_n722), .Y(
        aes_core_keymem_n2423) );
  AOI22X1 aes_core_keymem_U1541 ( .A0(aes_core_keymem_n2587), .A1(
        aes_core_keymem_n725), .B0(Din[172]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n724) );
  BUFX3 aes_core_keymem_U1540 ( .A(aes_core_keymem_n724), .Y(
        aes_core_keymem_n2422) );
  AOI22X1 aes_core_keymem_U1539 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n727), .B0(Din[171]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n726) );
  BUFX3 aes_core_keymem_U1538 ( .A(aes_core_keymem_n726), .Y(
        aes_core_keymem_n2421) );
  AOI22X1 aes_core_keymem_U1537 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n729), .B0(Din[170]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n728) );
  BUFX3 aes_core_keymem_U1536 ( .A(aes_core_keymem_n728), .Y(
        aes_core_keymem_n2420) );
  AOI22X1 aes_core_keymem_U1535 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n731), .B0(Din[169]), .B1(aes_core_keymem_n1), .Y(
        aes_core_keymem_n730) );
  BUFX3 aes_core_keymem_U1534 ( .A(aes_core_keymem_n730), .Y(
        aes_core_keymem_n2419) );
  AOI22X1 aes_core_keymem_U1533 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n733), .B0(Din[168]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n732) );
  BUFX3 aes_core_keymem_U1532 ( .A(aes_core_keymem_n732), .Y(
        aes_core_keymem_n2418) );
  AOI22X1 aes_core_keymem_U1531 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n735), .B0(Din[167]), .B1(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n734) );
  BUFX3 aes_core_keymem_U1530 ( .A(aes_core_keymem_n734), .Y(
        aes_core_keymem_n2417) );
  AOI22X1 aes_core_keymem_U1529 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n737), .B0(Din[166]), .B1(aes_core_keymem_n1), .Y(
        aes_core_keymem_n736) );
  BUFX3 aes_core_keymem_U1528 ( .A(aes_core_keymem_n736), .Y(
        aes_core_keymem_n2416) );
  AOI22X1 aes_core_keymem_U1527 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n739), .B0(Din[165]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n738) );
  BUFX3 aes_core_keymem_U1526 ( .A(aes_core_keymem_n738), .Y(
        aes_core_keymem_n2415) );
  AOI22X1 aes_core_keymem_U1525 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n741), .B0(Din[164]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n740) );
  BUFX3 aes_core_keymem_U1524 ( .A(aes_core_keymem_n740), .Y(
        aes_core_keymem_n2414) );
  AOI22X1 aes_core_keymem_U1523 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n743), .B0(Din[163]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n742) );
  BUFX3 aes_core_keymem_U1522 ( .A(aes_core_keymem_n742), .Y(
        aes_core_keymem_n2413) );
  AOI22X1 aes_core_keymem_U1521 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n745), .B0(Din[162]), .B1(aes_core_keymem_n1), .Y(
        aes_core_keymem_n744) );
  BUFX3 aes_core_keymem_U1520 ( .A(aes_core_keymem_n744), .Y(
        aes_core_keymem_n2412) );
  AOI22X1 aes_core_keymem_U1519 ( .A0(aes_core_keymem_n2588), .A1(
        aes_core_keymem_n749), .B0(Din[160]), .B1(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n748) );
  BUFX3 aes_core_keymem_U1518 ( .A(aes_core_keymem_n748), .Y(
        aes_core_keymem_n2410) );
  AOI22X1 aes_core_keymem_U1517 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n754), .B0(Din[158]), .B1(aes_core_keymem_n2525), .Y(
        aes_core_keymem_n753) );
  AOI22X1 aes_core_keymem_U1516 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n757), .B0(Din[157]), .B1(aes_core_keymem_n2551), .Y(
        aes_core_keymem_n756) );
  AOI22X1 aes_core_keymem_U1515 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n760), .B0(Din[156]), .B1(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n759) );
  AOI22X1 aes_core_keymem_U1514 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n763), .B0(Din[155]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n762) );
  AOI22X1 aes_core_keymem_U1513 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n772), .B0(Din[152]), .B1(aes_core_keymem_n2523), .Y(
        aes_core_keymem_n771) );
  AOI22X1 aes_core_keymem_U1512 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n775), .B0(Din[151]), .B1(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n774) );
  AOI22X1 aes_core_keymem_U1511 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n777), .B0(Din[150]), .B1(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n776) );
  AOI22X1 aes_core_keymem_U1510 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n779), .B0(Din[149]), .B1(aes_core_keymem_n2526), .Y(
        aes_core_keymem_n778) );
  AOI22X1 aes_core_keymem_U1509 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n781), .B0(Din[148]), .B1(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n780) );
  AOI22X1 aes_core_keymem_U1508 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n783), .B0(Din[147]), .B1(aes_core_keymem_n2525), .Y(
        aes_core_keymem_n782) );
  AOI22X1 aes_core_keymem_U1507 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n785), .B0(Din[146]), .B1(aes_core_keymem_n1), .Y(
        aes_core_keymem_n784) );
  AOI22X1 aes_core_keymem_U1506 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n787), .B0(Din[145]), .B1(aes_core_keymem_n2522), .Y(
        aes_core_keymem_n786) );
  AOI22X1 aes_core_keymem_U1505 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n789), .B0(Din[144]), .B1(aes_core_keymem_n2526), .Y(
        aes_core_keymem_n788) );
  AOI22X1 aes_core_keymem_U1504 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n793), .B0(Din[142]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n792) );
  AOI22X1 aes_core_keymem_U1503 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n795), .B0(Din[141]), .B1(aes_core_keymem_n2524), .Y(
        aes_core_keymem_n794) );
  AOI22X1 aes_core_keymem_U1502 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n797), .B0(Din[140]), .B1(aes_core_keymem_n2522), .Y(
        aes_core_keymem_n796) );
  AOI22X1 aes_core_keymem_U1501 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n799), .B0(Din[139]), .B1(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n798) );
  AOI22X1 aes_core_keymem_U1500 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n805), .B0(Din[136]), .B1(aes_core_keymem_n2552), .Y(
        aes_core_keymem_n804) );
  XOR2X1 aes_core_keymem_U1499 ( .A(aes_core_keymem_n737), .B(
        aes_core_keymem_sboxw[6]), .Y(aes_core_keymem_n809) );
  XOR2X1 aes_core_keymem_U1498 ( .A(aes_core_keymem_n739), .B(
        aes_core_keymem_sboxw[5]), .Y(aes_core_keymem_n811) );
  XOR2X1 aes_core_keymem_U1497 ( .A(aes_core_keymem_n741), .B(
        aes_core_keymem_sboxw[4]), .Y(aes_core_keymem_n813) );
  AOI22X1 aes_core_keymem_U1496 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n815), .B0(Din[131]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n814) );
  XOR2X1 aes_core_keymem_U1495 ( .A(aes_core_keymem_n745), .B(
        aes_core_keymem_sboxw[2]), .Y(aes_core_keymem_n817) );
  XOR2X1 aes_core_keymem_U1494 ( .A(aes_core_keymem_n747), .B(
        aes_core_keymem_sboxw[1]), .Y(aes_core_keymem_n819) );
  XOR2X1 aes_core_keymem_U1493 ( .A(aes_core_keymem_n749), .B(
        aes_core_keymem_sboxw[0]), .Y(aes_core_keymem_n830) );
  XOR2X1 aes_core_keymem_U1492 ( .A(aes_core_keymem_n625), .B(
        aes_core_keymem_prev_key1_reg[62]), .Y(aes_core_keymem_n689) );
  XOR2X1 aes_core_keymem_U1491 ( .A(aes_core_keymem_n627), .B(
        aes_core_keymem_prev_key1_reg[61]), .Y(aes_core_keymem_n691) );
  XOR2X1 aes_core_keymem_U1490 ( .A(aes_core_keymem_n629), .B(
        aes_core_keymem_prev_key1_reg[60]), .Y(aes_core_keymem_n693) );
  XOR2X1 aes_core_keymem_U1489 ( .A(aes_core_keymem_n631), .B(
        aes_core_keymem_prev_key1_reg[59]), .Y(aes_core_keymem_n695) );
  XOR2X1 aes_core_keymem_U1488 ( .A(aes_core_keymem_n633), .B(
        aes_core_keymem_prev_key1_reg[58]), .Y(aes_core_keymem_n697) );
  XOR2X1 aes_core_keymem_U1487 ( .A(aes_core_keymem_n635), .B(
        aes_core_keymem_prev_key1_reg[57]), .Y(aes_core_keymem_n699) );
  XOR2X1 aes_core_keymem_U1486 ( .A(aes_core_keymem_n637), .B(
        aes_core_keymem_prev_key1_reg[56]), .Y(aes_core_keymem_n701) );
  XOR2X1 aes_core_keymem_U1485 ( .A(aes_core_keymem_n639), .B(
        aes_core_keymem_prev_key1_reg[55]), .Y(aes_core_keymem_n703) );
  XOR2X1 aes_core_keymem_U1484 ( .A(aes_core_keymem_n641), .B(
        aes_core_keymem_prev_key1_reg[54]), .Y(aes_core_keymem_n705) );
  XOR2X1 aes_core_keymem_U1483 ( .A(aes_core_keymem_n643), .B(
        aes_core_keymem_prev_key1_reg[53]), .Y(aes_core_keymem_n707) );
  XOR2X1 aes_core_keymem_U1482 ( .A(aes_core_keymem_n645), .B(
        aes_core_keymem_prev_key1_reg[52]), .Y(aes_core_keymem_n709) );
  XOR2X1 aes_core_keymem_U1481 ( .A(aes_core_keymem_n647), .B(
        aes_core_keymem_prev_key1_reg[51]), .Y(aes_core_keymem_n711) );
  XOR2X1 aes_core_keymem_U1480 ( .A(aes_core_keymem_n649), .B(
        aes_core_keymem_prev_key1_reg[50]), .Y(aes_core_keymem_n713) );
  XOR2X1 aes_core_keymem_U1479 ( .A(aes_core_keymem_n651), .B(
        aes_core_keymem_prev_key1_reg[49]), .Y(aes_core_keymem_n715) );
  XOR2X1 aes_core_keymem_U1478 ( .A(aes_core_keymem_n653), .B(
        aes_core_keymem_prev_key1_reg[48]), .Y(aes_core_keymem_n717) );
  XOR2X1 aes_core_keymem_U1477 ( .A(aes_core_keymem_n657), .B(
        aes_core_keymem_prev_key1_reg[46]), .Y(aes_core_keymem_n721) );
  XOR2X1 aes_core_keymem_U1476 ( .A(aes_core_keymem_n659), .B(
        aes_core_keymem_prev_key1_reg[45]), .Y(aes_core_keymem_n723) );
  XOR2X1 aes_core_keymem_U1475 ( .A(aes_core_keymem_n661), .B(
        aes_core_keymem_prev_key1_reg[44]), .Y(aes_core_keymem_n725) );
  XOR2X1 aes_core_keymem_U1474 ( .A(aes_core_keymem_n663), .B(
        aes_core_keymem_prev_key1_reg[43]), .Y(aes_core_keymem_n727) );
  XOR2X1 aes_core_keymem_U1473 ( .A(aes_core_keymem_n665), .B(
        aes_core_keymem_prev_key1_reg[42]), .Y(aes_core_keymem_n729) );
  XOR2X1 aes_core_keymem_U1472 ( .A(aes_core_keymem_n667), .B(
        aes_core_keymem_prev_key1_reg[41]), .Y(aes_core_keymem_n731) );
  XOR2X1 aes_core_keymem_U1471 ( .A(aes_core_keymem_n669), .B(
        aes_core_keymem_prev_key1_reg[40]), .Y(aes_core_keymem_n733) );
  XOR2X1 aes_core_keymem_U1470 ( .A(aes_core_keymem_n671), .B(
        aes_core_keymem_prev_key1_reg[39]), .Y(aes_core_keymem_n735) );
  XOR2X1 aes_core_keymem_U1469 ( .A(aes_core_keymem_n673), .B(
        aes_core_keymem_prev_key1_reg[38]), .Y(aes_core_keymem_n737) );
  XOR2X1 aes_core_keymem_U1468 ( .A(aes_core_keymem_n675), .B(
        aes_core_keymem_prev_key1_reg[37]), .Y(aes_core_keymem_n739) );
  XOR2X1 aes_core_keymem_U1467 ( .A(aes_core_keymem_n677), .B(
        aes_core_keymem_prev_key1_reg[36]), .Y(aes_core_keymem_n741) );
  XOR2X1 aes_core_keymem_U1466 ( .A(aes_core_keymem_n679), .B(
        aes_core_keymem_prev_key1_reg[35]), .Y(aes_core_keymem_n743) );
  XOR2X1 aes_core_keymem_U1465 ( .A(aes_core_keymem_n681), .B(
        aes_core_keymem_prev_key1_reg[34]), .Y(aes_core_keymem_n745) );
  XOR2X1 aes_core_keymem_U1464 ( .A(aes_core_keymem_n683), .B(
        aes_core_keymem_prev_key1_reg[33]), .Y(aes_core_keymem_n747) );
  XOR2X1 aes_core_keymem_U1463 ( .A(aes_core_keymem_n685), .B(
        aes_core_keymem_prev_key1_reg[32]), .Y(aes_core_keymem_n749) );
  AOI22X1 aes_core_keymem_U1462 ( .A0(aes_core_keymem_n2586), .A1(
        aes_core_keymem_n687), .B0(Din[191]), .B1(aes_core_keymem_n2550), .Y(
        aes_core_keymem_n686) );
  BUFX3 aes_core_keymem_U1461 ( .A(aes_core_keymem_n686), .Y(
        aes_core_keymem_n2441) );
  AOI22X1 aes_core_keymem_U1460 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n751), .B0(Din[159]), .B1(aes_core_keymem_n2552), .Y(
        aes_core_keymem_n750) );
  AOI22X1 aes_core_keymem_U1459 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n791), .B0(Din[143]), .B1(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n790) );
  XOR2X1 aes_core_keymem_U1458 ( .A(aes_core_keymem_n623), .B(
        aes_core_keymem_prev_key1_reg[63]), .Y(aes_core_keymem_n687) );
  XOR2X1 aes_core_keymem_U1457 ( .A(aes_core_keymem_n655), .B(
        aes_core_keymem_prev_key1_reg[47]), .Y(aes_core_keymem_n719) );
  INVX2 aes_core_keymem_U1456 ( .A(aes_core_keymem_round_ctr_reg[0]), .Y(
        aes_core_keymem_n2767) );
  OAI2BB2X1 aes_core_keymem_U1455 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[127]), .Y(aes_core_keymem_n853) );
  OAI2BB2X1 aes_core_keymem_U1454 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[126]), .Y(aes_core_keymem_n865) );
  OAI2BB2X1 aes_core_keymem_U1453 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[125]), .Y(aes_core_keymem_n877) );
  OAI2BB2X1 aes_core_keymem_U1452 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[124]), .Y(aes_core_keymem_n889) );
  OAI2BB2X1 aes_core_keymem_U1451 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[123]), .Y(aes_core_keymem_n901) );
  OAI2BB2X1 aes_core_keymem_U1450 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[122]), .Y(aes_core_keymem_n913) );
  OAI2BB2X1 aes_core_keymem_U1449 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[121]), .Y(aes_core_keymem_n925) );
  OAI2BB2X1 aes_core_keymem_U1448 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[120]), .Y(aes_core_keymem_n937) );
  OAI2BB2X1 aes_core_keymem_U1447 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[119]), .Y(aes_core_keymem_n949) );
  OAI2BB2X1 aes_core_keymem_U1446 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[118]), .Y(aes_core_keymem_n961) );
  OAI2BB2X1 aes_core_keymem_U1445 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[117]), .Y(aes_core_keymem_n973) );
  OAI2BB2X1 aes_core_keymem_U1444 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[116]), .Y(aes_core_keymem_n985) );
  OAI2BB2X1 aes_core_keymem_U1443 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[115]), .Y(aes_core_keymem_n997) );
  OAI2BB2X1 aes_core_keymem_U1442 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[114]), .Y(aes_core_keymem_n1009) );
  OAI2BB2X1 aes_core_keymem_U1441 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[113]), .Y(aes_core_keymem_n1021) );
  OAI2BB2X1 aes_core_keymem_U1440 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[112]), .Y(aes_core_keymem_n1033) );
  OAI2BB2X1 aes_core_keymem_U1439 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[111]), .Y(aes_core_keymem_n1045) );
  OAI2BB2X1 aes_core_keymem_U1438 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[110]), .Y(aes_core_keymem_n1057) );
  OAI2BB2X1 aes_core_keymem_U1437 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[109]), .Y(aes_core_keymem_n1069) );
  OAI2BB2X1 aes_core_keymem_U1436 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[108]), .Y(aes_core_keymem_n1081) );
  OAI2BB2X1 aes_core_keymem_U1435 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[107]), .Y(aes_core_keymem_n1093) );
  OAI2BB2X1 aes_core_keymem_U1434 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[106]), .Y(aes_core_keymem_n1105) );
  OAI2BB2X1 aes_core_keymem_U1433 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[105]), .Y(aes_core_keymem_n1117) );
  OAI2BB2X1 aes_core_keymem_U1432 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[104]), .Y(aes_core_keymem_n1129) );
  OAI2BB2X1 aes_core_keymem_U1431 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[103]), .Y(aes_core_keymem_n1141) );
  OAI2BB2X1 aes_core_keymem_U1430 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[102]), .Y(aes_core_keymem_n1153) );
  OAI2BB2X1 aes_core_keymem_U1429 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[101]), .Y(aes_core_keymem_n1165) );
  OAI2BB2X1 aes_core_keymem_U1428 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[100]), .Y(aes_core_keymem_n1177) );
  OAI2BB2X1 aes_core_keymem_U1427 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[99]), .Y(aes_core_keymem_n1189) );
  OAI2BB2X1 aes_core_keymem_U1426 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[98]), .Y(aes_core_keymem_n1201) );
  OAI2BB2X1 aes_core_keymem_U1425 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[97]), .Y(aes_core_keymem_n1213) );
  OAI2BB2X1 aes_core_keymem_U1424 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[96]), .Y(aes_core_keymem_n1225) );
  OAI2BB2X1 aes_core_keymem_U1423 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[95]), .Y(aes_core_keymem_n1237) );
  OAI2BB2X1 aes_core_keymem_U1422 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[94]), .Y(aes_core_keymem_n1249) );
  OAI2BB2X1 aes_core_keymem_U1421 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[93]), .Y(aes_core_keymem_n1261) );
  OAI2BB2X1 aes_core_keymem_U1420 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[92]), .Y(aes_core_keymem_n1273) );
  OAI2BB2X1 aes_core_keymem_U1419 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[91]), .Y(aes_core_keymem_n1285) );
  OAI2BB2X1 aes_core_keymem_U1418 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[90]), .Y(aes_core_keymem_n1297) );
  OAI2BB2X1 aes_core_keymem_U1417 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[89]), .Y(aes_core_keymem_n1309) );
  OAI2BB2X1 aes_core_keymem_U1416 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[88]), .Y(aes_core_keymem_n1321) );
  OAI2BB2X1 aes_core_keymem_U1415 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[87]), .Y(aes_core_keymem_n1333) );
  OAI2BB2X1 aes_core_keymem_U1414 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[86]), .Y(aes_core_keymem_n1345) );
  OAI2BB2X1 aes_core_keymem_U1413 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[85]), .Y(aes_core_keymem_n1357) );
  OAI2BB2X1 aes_core_keymem_U1412 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[84]), .Y(aes_core_keymem_n1369) );
  OAI2BB2X1 aes_core_keymem_U1411 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[83]), .Y(aes_core_keymem_n1381) );
  OAI2BB2X1 aes_core_keymem_U1410 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[82]), .Y(aes_core_keymem_n1393) );
  OAI2BB2X1 aes_core_keymem_U1409 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[81]), .Y(aes_core_keymem_n1405) );
  OAI2BB2X1 aes_core_keymem_U1408 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[80]), .Y(aes_core_keymem_n1417) );
  OAI2BB2X1 aes_core_keymem_U1407 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[79]), .Y(aes_core_keymem_n1429) );
  OAI2BB2X1 aes_core_keymem_U1406 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[78]), .Y(aes_core_keymem_n1441) );
  OAI2BB2X1 aes_core_keymem_U1405 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[77]), .Y(aes_core_keymem_n1453) );
  OAI2BB2X1 aes_core_keymem_U1404 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[76]), .Y(aes_core_keymem_n1465) );
  OAI2BB2X1 aes_core_keymem_U1403 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[75]), .Y(aes_core_keymem_n1477) );
  OAI2BB2X1 aes_core_keymem_U1402 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[74]), .Y(aes_core_keymem_n1489) );
  OAI2BB2X1 aes_core_keymem_U1401 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[73]), .Y(aes_core_keymem_n1501) );
  OAI2BB2X1 aes_core_keymem_U1400 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[72]), .Y(aes_core_keymem_n1513) );
  OAI2BB2X1 aes_core_keymem_U1399 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[71]), .Y(aes_core_keymem_n1525) );
  OAI2BB2X1 aes_core_keymem_U1398 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[70]), .Y(aes_core_keymem_n1537) );
  OAI2BB2X1 aes_core_keymem_U1397 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[69]), .Y(aes_core_keymem_n1549) );
  OAI2BB2X1 aes_core_keymem_U1396 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[68]), .Y(aes_core_keymem_n1561) );
  OAI2BB2X1 aes_core_keymem_U1395 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[67]), .Y(aes_core_keymem_n1573) );
  OAI2BB2X1 aes_core_keymem_U1394 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[66]), .Y(aes_core_keymem_n1585) );
  OAI2BB2X1 aes_core_keymem_U1393 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[65]), .Y(aes_core_keymem_n1597) );
  OAI2BB2X1 aes_core_keymem_U1392 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[64]), .Y(aes_core_keymem_n1609) );
  OAI2BB2X1 aes_core_keymem_U1391 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[63]), .Y(aes_core_keymem_n1621) );
  OAI2BB2X1 aes_core_keymem_U1390 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[62]), .Y(aes_core_keymem_n1633) );
  OAI2BB2X1 aes_core_keymem_U1389 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[61]), .Y(aes_core_keymem_n1645) );
  OAI2BB2X1 aes_core_keymem_U1388 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[60]), .Y(aes_core_keymem_n1657) );
  OAI2BB2X1 aes_core_keymem_U1387 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[59]), .Y(aes_core_keymem_n1669) );
  OAI2BB2X1 aes_core_keymem_U1386 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[58]), .Y(aes_core_keymem_n1681) );
  OAI2BB2X1 aes_core_keymem_U1385 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[57]), .Y(aes_core_keymem_n1693) );
  OAI2BB2X1 aes_core_keymem_U1384 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[56]), .Y(aes_core_keymem_n1705) );
  OAI2BB2X1 aes_core_keymem_U1383 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[55]), .Y(aes_core_keymem_n1717) );
  OAI2BB2X1 aes_core_keymem_U1382 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[54]), .Y(aes_core_keymem_n1729) );
  OAI2BB2X1 aes_core_keymem_U1381 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[53]), .Y(aes_core_keymem_n1741) );
  OAI2BB2X1 aes_core_keymem_U1380 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[52]), .Y(aes_core_keymem_n1753) );
  OAI2BB2X1 aes_core_keymem_U1379 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[51]), .Y(aes_core_keymem_n1765) );
  OAI2BB2X1 aes_core_keymem_U1378 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[50]), .Y(aes_core_keymem_n1777) );
  OAI2BB2X1 aes_core_keymem_U1377 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[49]), .Y(aes_core_keymem_n1789) );
  OAI2BB2X1 aes_core_keymem_U1376 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[48]), .Y(aes_core_keymem_n1801) );
  OAI2BB2X1 aes_core_keymem_U1375 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[47]), .Y(aes_core_keymem_n1813) );
  OAI2BB2X1 aes_core_keymem_U1374 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[46]), .Y(aes_core_keymem_n1825) );
  OAI2BB2X1 aes_core_keymem_U1373 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[45]), .Y(aes_core_keymem_n1837) );
  OAI2BB2X1 aes_core_keymem_U1372 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[44]), .Y(aes_core_keymem_n1849) );
  OAI2BB2X1 aes_core_keymem_U1371 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[43]), .Y(aes_core_keymem_n1861) );
  OAI2BB2X1 aes_core_keymem_U1370 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[42]), .Y(aes_core_keymem_n1873) );
  OAI2BB2X1 aes_core_keymem_U1369 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[41]), .Y(aes_core_keymem_n1885) );
  OAI2BB2X1 aes_core_keymem_U1368 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[40]), .Y(aes_core_keymem_n1897) );
  OAI2BB2X1 aes_core_keymem_U1367 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[39]), .Y(aes_core_keymem_n1909) );
  OAI2BB2X1 aes_core_keymem_U1366 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[38]), .Y(aes_core_keymem_n1921) );
  OAI2BB2X1 aes_core_keymem_U1365 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[37]), .Y(aes_core_keymem_n1933) );
  OAI2BB2X1 aes_core_keymem_U1364 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[36]), .Y(aes_core_keymem_n1945) );
  OAI2BB2X1 aes_core_keymem_U1363 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[35]), .Y(aes_core_keymem_n1957) );
  OAI2BB2X1 aes_core_keymem_U1362 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[34]), .Y(aes_core_keymem_n1969) );
  OAI2BB2X1 aes_core_keymem_U1361 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[33]), .Y(aes_core_keymem_n1981) );
  OAI2BB2X1 aes_core_keymem_U1360 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_prev_key1_reg[32]), .Y(aes_core_keymem_n1993) );
  OAI2BB2X1 aes_core_keymem_U1359 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[31]), .Y(aes_core_keymem_n2005) );
  OAI2BB2X1 aes_core_keymem_U1358 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[30]), .Y(aes_core_keymem_n2017) );
  OAI2BB2X1 aes_core_keymem_U1357 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[29]), .Y(aes_core_keymem_n2029) );
  OAI2BB2X1 aes_core_keymem_U1356 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[28]), .Y(aes_core_keymem_n2041) );
  OAI2BB2X1 aes_core_keymem_U1355 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[27]), .Y(aes_core_keymem_n2053) );
  OAI2BB2X1 aes_core_keymem_U1354 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[26]), .Y(aes_core_keymem_n2065) );
  OAI2BB2X1 aes_core_keymem_U1353 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[25]), .Y(aes_core_keymem_n2077) );
  OAI2BB2X1 aes_core_keymem_U1352 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[24]), .Y(aes_core_keymem_n2089) );
  OAI2BB2X1 aes_core_keymem_U1351 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[23]), .Y(aes_core_keymem_n2101) );
  OAI2BB2X1 aes_core_keymem_U1350 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[22]), .Y(aes_core_keymem_n2113) );
  OAI2BB2X1 aes_core_keymem_U1349 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[21]), .Y(aes_core_keymem_n2125) );
  OAI2BB2X1 aes_core_keymem_U1348 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[20]), .Y(aes_core_keymem_n2137) );
  OAI2BB2X1 aes_core_keymem_U1347 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[19]), .Y(aes_core_keymem_n2149) );
  OAI2BB2X1 aes_core_keymem_U1346 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[18]), .Y(aes_core_keymem_n2161) );
  OAI2BB2X1 aes_core_keymem_U1345 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[17]), .Y(aes_core_keymem_n2173) );
  OAI2BB2X1 aes_core_keymem_U1344 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[16]), .Y(aes_core_keymem_n2185) );
  OAI2BB2X1 aes_core_keymem_U1343 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[15]), .Y(aes_core_keymem_n2197) );
  OAI2BB2X1 aes_core_keymem_U1342 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[14]), .Y(aes_core_keymem_n2209) );
  OAI2BB2X1 aes_core_keymem_U1341 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[13]), .Y(aes_core_keymem_n2221) );
  OAI2BB2X1 aes_core_keymem_U1340 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[12]), .Y(aes_core_keymem_n2233) );
  OAI2BB2X1 aes_core_keymem_U1339 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[11]), .Y(aes_core_keymem_n2245) );
  OAI2BB2X1 aes_core_keymem_U1338 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[10]), .Y(aes_core_keymem_n2257) );
  OAI2BB2X1 aes_core_keymem_U1337 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[9]), .Y(aes_core_keymem_n2269) );
  OAI2BB2X1 aes_core_keymem_U1336 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[8]), .Y(aes_core_keymem_n2281) );
  OAI2BB2X1 aes_core_keymem_U1335 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[7]), .Y(aes_core_keymem_n2293) );
  OAI2BB2X1 aes_core_keymem_U1334 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[6]), .Y(aes_core_keymem_n2305) );
  OAI2BB2X1 aes_core_keymem_U1333 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[5]), .Y(aes_core_keymem_n2317) );
  OAI2BB2X1 aes_core_keymem_U1332 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[4]), .Y(aes_core_keymem_n2329) );
  OAI2BB2X1 aes_core_keymem_U1331 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[3]), .Y(aes_core_keymem_n2341) );
  OAI2BB2X1 aes_core_keymem_U1330 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[2]), .Y(aes_core_keymem_n2353) );
  OAI2BB2X1 aes_core_keymem_U1329 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[1]), .Y(aes_core_keymem_n2365) );
  OAI2BB2X1 aes_core_keymem_U1328 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n9), .A0N(aes_core_keymem_n9), .A1N(
        aes_core_keymem_sboxw[0]), .Y(aes_core_keymem_n2377) );
  OAI2BB2X1 aes_core_keymem_U1327 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[895]), .Y(aes_core_keymem_n844) );
  OAI2BB2X1 aes_core_keymem_U1326 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[894]), .Y(aes_core_keymem_n856) );
  OAI2BB2X1 aes_core_keymem_U1325 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[893]), .Y(aes_core_keymem_n868) );
  OAI2BB2X1 aes_core_keymem_U1324 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[892]), .Y(aes_core_keymem_n880) );
  OAI2BB2X1 aes_core_keymem_U1323 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[891]), .Y(aes_core_keymem_n892) );
  OAI2BB2X1 aes_core_keymem_U1322 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[890]), .Y(aes_core_keymem_n904) );
  OAI2BB2X1 aes_core_keymem_U1321 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[889]), .Y(aes_core_keymem_n916) );
  OAI2BB2X1 aes_core_keymem_U1320 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[888]), .Y(aes_core_keymem_n928) );
  OAI2BB2X1 aes_core_keymem_U1319 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[887]), .Y(aes_core_keymem_n940) );
  OAI2BB2X1 aes_core_keymem_U1318 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[886]), .Y(aes_core_keymem_n952) );
  OAI2BB2X1 aes_core_keymem_U1317 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[885]), .Y(aes_core_keymem_n964) );
  OAI2BB2X1 aes_core_keymem_U1316 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[884]), .Y(aes_core_keymem_n976) );
  OAI2BB2X1 aes_core_keymem_U1315 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[883]), .Y(aes_core_keymem_n988) );
  OAI2BB2X1 aes_core_keymem_U1314 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[882]), .Y(aes_core_keymem_n1000) );
  OAI2BB2X1 aes_core_keymem_U1313 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[881]), .Y(aes_core_keymem_n1012) );
  OAI2BB2X1 aes_core_keymem_U1312 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[880]), .Y(aes_core_keymem_n1024) );
  OAI2BB2X1 aes_core_keymem_U1311 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[879]), .Y(aes_core_keymem_n1036) );
  OAI2BB2X1 aes_core_keymem_U1310 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[878]), .Y(aes_core_keymem_n1048) );
  OAI2BB2X1 aes_core_keymem_U1309 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[877]), .Y(aes_core_keymem_n1060) );
  OAI2BB2X1 aes_core_keymem_U1308 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[876]), .Y(aes_core_keymem_n1072) );
  OAI2BB2X1 aes_core_keymem_U1307 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[875]), .Y(aes_core_keymem_n1084) );
  OAI2BB2X1 aes_core_keymem_U1306 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[874]), .Y(aes_core_keymem_n1096) );
  OAI2BB2X1 aes_core_keymem_U1305 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[873]), .Y(aes_core_keymem_n1108) );
  OAI2BB2X1 aes_core_keymem_U1304 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[872]), .Y(aes_core_keymem_n1120) );
  OAI2BB2X1 aes_core_keymem_U1303 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[871]), .Y(aes_core_keymem_n1132) );
  OAI2BB2X1 aes_core_keymem_U1302 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[870]), .Y(aes_core_keymem_n1144) );
  OAI2BB2X1 aes_core_keymem_U1301 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[869]), .Y(aes_core_keymem_n1156) );
  OAI2BB2X1 aes_core_keymem_U1300 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[868]), .Y(aes_core_keymem_n1168) );
  OAI2BB2X1 aes_core_keymem_U1299 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[867]), .Y(aes_core_keymem_n1180) );
  OAI2BB2X1 aes_core_keymem_U1298 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[866]), .Y(aes_core_keymem_n1192) );
  OAI2BB2X1 aes_core_keymem_U1297 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[865]), .Y(aes_core_keymem_n1204) );
  OAI2BB2X1 aes_core_keymem_U1296 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[864]), .Y(aes_core_keymem_n1216) );
  OAI2BB2X1 aes_core_keymem_U1295 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[863]), .Y(aes_core_keymem_n1228) );
  OAI2BB2X1 aes_core_keymem_U1294 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[862]), .Y(aes_core_keymem_n1240) );
  OAI2BB2X1 aes_core_keymem_U1293 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[861]), .Y(aes_core_keymem_n1252) );
  OAI2BB2X1 aes_core_keymem_U1292 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[860]), .Y(aes_core_keymem_n1264) );
  OAI2BB2X1 aes_core_keymem_U1291 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[859]), .Y(aes_core_keymem_n1276) );
  OAI2BB2X1 aes_core_keymem_U1290 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[858]), .Y(aes_core_keymem_n1288) );
  OAI2BB2X1 aes_core_keymem_U1289 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[857]), .Y(aes_core_keymem_n1300) );
  OAI2BB2X1 aes_core_keymem_U1288 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[856]), .Y(aes_core_keymem_n1312) );
  OAI2BB2X1 aes_core_keymem_U1287 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[855]), .Y(aes_core_keymem_n1324) );
  OAI2BB2X1 aes_core_keymem_U1286 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[854]), .Y(aes_core_keymem_n1336) );
  OAI2BB2X1 aes_core_keymem_U1285 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[853]), .Y(aes_core_keymem_n1348) );
  OAI2BB2X1 aes_core_keymem_U1284 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[852]), .Y(aes_core_keymem_n1360) );
  OAI2BB2X1 aes_core_keymem_U1283 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[851]), .Y(aes_core_keymem_n1372) );
  OAI2BB2X1 aes_core_keymem_U1282 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[850]), .Y(aes_core_keymem_n1384) );
  OAI2BB2X1 aes_core_keymem_U1281 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[849]), .Y(aes_core_keymem_n1396) );
  OAI2BB2X1 aes_core_keymem_U1280 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[848]), .Y(aes_core_keymem_n1408) );
  OAI2BB2X1 aes_core_keymem_U1279 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[847]), .Y(aes_core_keymem_n1420) );
  OAI2BB2X1 aes_core_keymem_U1278 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[846]), .Y(aes_core_keymem_n1432) );
  OAI2BB2X1 aes_core_keymem_U1277 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[845]), .Y(aes_core_keymem_n1444) );
  OAI2BB2X1 aes_core_keymem_U1276 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[844]), .Y(aes_core_keymem_n1456) );
  OAI2BB2X1 aes_core_keymem_U1275 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[843]), .Y(aes_core_keymem_n1468) );
  OAI2BB2X1 aes_core_keymem_U1274 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[842]), .Y(aes_core_keymem_n1480) );
  OAI2BB2X1 aes_core_keymem_U1273 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[841]), .Y(aes_core_keymem_n1492) );
  OAI2BB2X1 aes_core_keymem_U1272 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[840]), .Y(aes_core_keymem_n1504) );
  OAI2BB2X1 aes_core_keymem_U1271 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[839]), .Y(aes_core_keymem_n1516) );
  OAI2BB2X1 aes_core_keymem_U1270 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[838]), .Y(aes_core_keymem_n1528) );
  OAI2BB2X1 aes_core_keymem_U1269 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[837]), .Y(aes_core_keymem_n1540) );
  OAI2BB2X1 aes_core_keymem_U1268 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[836]), .Y(aes_core_keymem_n1552) );
  OAI2BB2X1 aes_core_keymem_U1267 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[835]), .Y(aes_core_keymem_n1564) );
  OAI2BB2X1 aes_core_keymem_U1266 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[834]), .Y(aes_core_keymem_n1576) );
  OAI2BB2X1 aes_core_keymem_U1265 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[833]), .Y(aes_core_keymem_n1588) );
  OAI2BB2X1 aes_core_keymem_U1264 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[832]), .Y(aes_core_keymem_n1600) );
  OAI2BB2X1 aes_core_keymem_U1263 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[831]), .Y(aes_core_keymem_n1612) );
  OAI2BB2X1 aes_core_keymem_U1262 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[830]), .Y(aes_core_keymem_n1624) );
  OAI2BB2X1 aes_core_keymem_U1261 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[829]), .Y(aes_core_keymem_n1636) );
  OAI2BB2X1 aes_core_keymem_U1260 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[828]), .Y(aes_core_keymem_n1648) );
  OAI2BB2X1 aes_core_keymem_U1259 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[827]), .Y(aes_core_keymem_n1660) );
  OAI2BB2X1 aes_core_keymem_U1258 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[826]), .Y(aes_core_keymem_n1672) );
  OAI2BB2X1 aes_core_keymem_U1257 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[825]), .Y(aes_core_keymem_n1684) );
  OAI2BB2X1 aes_core_keymem_U1256 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[824]), .Y(aes_core_keymem_n1696) );
  OAI2BB2X1 aes_core_keymem_U1255 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[823]), .Y(aes_core_keymem_n1708) );
  OAI2BB2X1 aes_core_keymem_U1254 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[822]), .Y(aes_core_keymem_n1720) );
  OAI2BB2X1 aes_core_keymem_U1253 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[821]), .Y(aes_core_keymem_n1732) );
  OAI2BB2X1 aes_core_keymem_U1252 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[820]), .Y(aes_core_keymem_n1744) );
  OAI2BB2X1 aes_core_keymem_U1251 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[819]), .Y(aes_core_keymem_n1756) );
  OAI2BB2X1 aes_core_keymem_U1250 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[818]), .Y(aes_core_keymem_n1768) );
  OAI2BB2X1 aes_core_keymem_U1249 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[817]), .Y(aes_core_keymem_n1780) );
  OAI2BB2X1 aes_core_keymem_U1248 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[816]), .Y(aes_core_keymem_n1792) );
  OAI2BB2X1 aes_core_keymem_U1247 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[815]), .Y(aes_core_keymem_n1804) );
  OAI2BB2X1 aes_core_keymem_U1246 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[814]), .Y(aes_core_keymem_n1816) );
  OAI2BB2X1 aes_core_keymem_U1245 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[813]), .Y(aes_core_keymem_n1828) );
  OAI2BB2X1 aes_core_keymem_U1244 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[812]), .Y(aes_core_keymem_n1840) );
  OAI2BB2X1 aes_core_keymem_U1243 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[811]), .Y(aes_core_keymem_n1852) );
  OAI2BB2X1 aes_core_keymem_U1242 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[810]), .Y(aes_core_keymem_n1864) );
  OAI2BB2X1 aes_core_keymem_U1241 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[809]), .Y(aes_core_keymem_n1876) );
  OAI2BB2X1 aes_core_keymem_U1240 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[808]), .Y(aes_core_keymem_n1888) );
  OAI2BB2X1 aes_core_keymem_U1239 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[807]), .Y(aes_core_keymem_n1900) );
  OAI2BB2X1 aes_core_keymem_U1238 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[806]), .Y(aes_core_keymem_n1912) );
  OAI2BB2X1 aes_core_keymem_U1237 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[805]), .Y(aes_core_keymem_n1924) );
  OAI2BB2X1 aes_core_keymem_U1236 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[804]), .Y(aes_core_keymem_n1936) );
  OAI2BB2X1 aes_core_keymem_U1235 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[803]), .Y(aes_core_keymem_n1948) );
  OAI2BB2X1 aes_core_keymem_U1234 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[802]), .Y(aes_core_keymem_n1960) );
  OAI2BB2X1 aes_core_keymem_U1233 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[801]), .Y(aes_core_keymem_n1972) );
  OAI2BB2X1 aes_core_keymem_U1232 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[800]), .Y(aes_core_keymem_n1984) );
  OAI2BB2X1 aes_core_keymem_U1231 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[799]), .Y(aes_core_keymem_n1996) );
  OAI2BB2X1 aes_core_keymem_U1230 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[798]), .Y(aes_core_keymem_n2008) );
  OAI2BB2X1 aes_core_keymem_U1229 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[797]), .Y(aes_core_keymem_n2020) );
  OAI2BB2X1 aes_core_keymem_U1228 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[796]), .Y(aes_core_keymem_n2032) );
  OAI2BB2X1 aes_core_keymem_U1227 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[795]), .Y(aes_core_keymem_n2044) );
  OAI2BB2X1 aes_core_keymem_U1226 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[794]), .Y(aes_core_keymem_n2056) );
  OAI2BB2X1 aes_core_keymem_U1225 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[793]), .Y(aes_core_keymem_n2068) );
  OAI2BB2X1 aes_core_keymem_U1224 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[792]), .Y(aes_core_keymem_n2080) );
  OAI2BB2X1 aes_core_keymem_U1223 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[791]), .Y(aes_core_keymem_n2092) );
  OAI2BB2X1 aes_core_keymem_U1222 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[790]), .Y(aes_core_keymem_n2104) );
  OAI2BB2X1 aes_core_keymem_U1221 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[789]), .Y(aes_core_keymem_n2116) );
  OAI2BB2X1 aes_core_keymem_U1220 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[788]), .Y(aes_core_keymem_n2128) );
  OAI2BB2X1 aes_core_keymem_U1219 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[787]), .Y(aes_core_keymem_n2140) );
  OAI2BB2X1 aes_core_keymem_U1218 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[786]), .Y(aes_core_keymem_n2152) );
  OAI2BB2X1 aes_core_keymem_U1217 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[785]), .Y(aes_core_keymem_n2164) );
  OAI2BB2X1 aes_core_keymem_U1216 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[784]), .Y(aes_core_keymem_n2176) );
  OAI2BB2X1 aes_core_keymem_U1215 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[783]), .Y(aes_core_keymem_n2188) );
  OAI2BB2X1 aes_core_keymem_U1214 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[782]), .Y(aes_core_keymem_n2200) );
  OAI2BB2X1 aes_core_keymem_U1213 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[781]), .Y(aes_core_keymem_n2212) );
  OAI2BB2X1 aes_core_keymem_U1212 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[780]), .Y(aes_core_keymem_n2224) );
  OAI2BB2X1 aes_core_keymem_U1211 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[779]), .Y(aes_core_keymem_n2236) );
  OAI2BB2X1 aes_core_keymem_U1210 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[778]), .Y(aes_core_keymem_n2248) );
  OAI2BB2X1 aes_core_keymem_U1209 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[777]), .Y(aes_core_keymem_n2260) );
  OAI2BB2X1 aes_core_keymem_U1208 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[776]), .Y(aes_core_keymem_n2272) );
  OAI2BB2X1 aes_core_keymem_U1207 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[775]), .Y(aes_core_keymem_n2284) );
  OAI2BB2X1 aes_core_keymem_U1206 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[774]), .Y(aes_core_keymem_n2296) );
  OAI2BB2X1 aes_core_keymem_U1205 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[773]), .Y(aes_core_keymem_n2308) );
  OAI2BB2X1 aes_core_keymem_U1204 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[772]), .Y(aes_core_keymem_n2320) );
  OAI2BB2X1 aes_core_keymem_U1203 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[771]), .Y(aes_core_keymem_n2332) );
  OAI2BB2X1 aes_core_keymem_U1202 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[770]), .Y(aes_core_keymem_n2344) );
  OAI2BB2X1 aes_core_keymem_U1201 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[769]), .Y(aes_core_keymem_n2356) );
  OAI2BB2X1 aes_core_keymem_U1200 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n549), .A0N(aes_core_keymem_n549), .A1N(
        aes_core_keymem_key_mem[768]), .Y(aes_core_keymem_n2368) );
  OAI2BB2X1 aes_core_keymem_U1199 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[767]), .Y(aes_core_keymem_n843) );
  OAI2BB2X1 aes_core_keymem_U1198 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[766]), .Y(aes_core_keymem_n855) );
  OAI2BB2X1 aes_core_keymem_U1197 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[765]), .Y(aes_core_keymem_n867) );
  OAI2BB2X1 aes_core_keymem_U1196 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[764]), .Y(aes_core_keymem_n879) );
  OAI2BB2X1 aes_core_keymem_U1195 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[763]), .Y(aes_core_keymem_n891) );
  OAI2BB2X1 aes_core_keymem_U1194 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[762]), .Y(aes_core_keymem_n903) );
  OAI2BB2X1 aes_core_keymem_U1193 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[761]), .Y(aes_core_keymem_n915) );
  OAI2BB2X1 aes_core_keymem_U1192 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[760]), .Y(aes_core_keymem_n927) );
  OAI2BB2X1 aes_core_keymem_U1191 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[759]), .Y(aes_core_keymem_n939) );
  OAI2BB2X1 aes_core_keymem_U1190 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[758]), .Y(aes_core_keymem_n951) );
  OAI2BB2X1 aes_core_keymem_U1189 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[757]), .Y(aes_core_keymem_n963) );
  OAI2BB2X1 aes_core_keymem_U1188 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[756]), .Y(aes_core_keymem_n975) );
  OAI2BB2X1 aes_core_keymem_U1187 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[755]), .Y(aes_core_keymem_n987) );
  OAI2BB2X1 aes_core_keymem_U1186 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[754]), .Y(aes_core_keymem_n999) );
  OAI2BB2X1 aes_core_keymem_U1185 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[753]), .Y(aes_core_keymem_n1011) );
  OAI2BB2X1 aes_core_keymem_U1184 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[752]), .Y(aes_core_keymem_n1023) );
  OAI2BB2X1 aes_core_keymem_U1183 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[751]), .Y(aes_core_keymem_n1035) );
  OAI2BB2X1 aes_core_keymem_U1182 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[750]), .Y(aes_core_keymem_n1047) );
  OAI2BB2X1 aes_core_keymem_U1181 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[749]), .Y(aes_core_keymem_n1059) );
  OAI2BB2X1 aes_core_keymem_U1180 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[748]), .Y(aes_core_keymem_n1071) );
  OAI2BB2X1 aes_core_keymem_U1179 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[747]), .Y(aes_core_keymem_n1083) );
  OAI2BB2X1 aes_core_keymem_U1178 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[746]), .Y(aes_core_keymem_n1095) );
  OAI2BB2X1 aes_core_keymem_U1177 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[745]), .Y(aes_core_keymem_n1107) );
  OAI2BB2X1 aes_core_keymem_U1176 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[744]), .Y(aes_core_keymem_n1119) );
  OAI2BB2X1 aes_core_keymem_U1175 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[743]), .Y(aes_core_keymem_n1131) );
  OAI2BB2X1 aes_core_keymem_U1174 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[742]), .Y(aes_core_keymem_n1143) );
  OAI2BB2X1 aes_core_keymem_U1173 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[741]), .Y(aes_core_keymem_n1155) );
  OAI2BB2X1 aes_core_keymem_U1172 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[740]), .Y(aes_core_keymem_n1167) );
  OAI2BB2X1 aes_core_keymem_U1171 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[739]), .Y(aes_core_keymem_n1179) );
  OAI2BB2X1 aes_core_keymem_U1170 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[738]), .Y(aes_core_keymem_n1191) );
  OAI2BB2X1 aes_core_keymem_U1169 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[737]), .Y(aes_core_keymem_n1203) );
  OAI2BB2X1 aes_core_keymem_U1168 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[736]), .Y(aes_core_keymem_n1215) );
  OAI2BB2X1 aes_core_keymem_U1167 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[735]), .Y(aes_core_keymem_n1227) );
  OAI2BB2X1 aes_core_keymem_U1166 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[734]), .Y(aes_core_keymem_n1239) );
  OAI2BB2X1 aes_core_keymem_U1165 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[733]), .Y(aes_core_keymem_n1251) );
  OAI2BB2X1 aes_core_keymem_U1164 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[732]), .Y(aes_core_keymem_n1263) );
  OAI2BB2X1 aes_core_keymem_U1163 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[731]), .Y(aes_core_keymem_n1275) );
  OAI2BB2X1 aes_core_keymem_U1162 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[730]), .Y(aes_core_keymem_n1287) );
  OAI2BB2X1 aes_core_keymem_U1161 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[729]), .Y(aes_core_keymem_n1299) );
  OAI2BB2X1 aes_core_keymem_U1160 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[728]), .Y(aes_core_keymem_n1311) );
  OAI2BB2X1 aes_core_keymem_U1159 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[727]), .Y(aes_core_keymem_n1323) );
  OAI2BB2X1 aes_core_keymem_U1158 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[726]), .Y(aes_core_keymem_n1335) );
  OAI2BB2X1 aes_core_keymem_U1157 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[725]), .Y(aes_core_keymem_n1347) );
  OAI2BB2X1 aes_core_keymem_U1156 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[724]), .Y(aes_core_keymem_n1359) );
  OAI2BB2X1 aes_core_keymem_U1155 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[723]), .Y(aes_core_keymem_n1371) );
  OAI2BB2X1 aes_core_keymem_U1154 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[722]), .Y(aes_core_keymem_n1383) );
  OAI2BB2X1 aes_core_keymem_U1153 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[721]), .Y(aes_core_keymem_n1395) );
  OAI2BB2X1 aes_core_keymem_U1152 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[720]), .Y(aes_core_keymem_n1407) );
  OAI2BB2X1 aes_core_keymem_U1151 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[719]), .Y(aes_core_keymem_n1419) );
  OAI2BB2X1 aes_core_keymem_U1150 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[718]), .Y(aes_core_keymem_n1431) );
  OAI2BB2X1 aes_core_keymem_U1149 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[717]), .Y(aes_core_keymem_n1443) );
  OAI2BB2X1 aes_core_keymem_U1148 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[716]), .Y(aes_core_keymem_n1455) );
  OAI2BB2X1 aes_core_keymem_U1147 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[715]), .Y(aes_core_keymem_n1467) );
  OAI2BB2X1 aes_core_keymem_U1146 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[714]), .Y(aes_core_keymem_n1479) );
  OAI2BB2X1 aes_core_keymem_U1145 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[713]), .Y(aes_core_keymem_n1491) );
  OAI2BB2X1 aes_core_keymem_U1144 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[712]), .Y(aes_core_keymem_n1503) );
  OAI2BB2X1 aes_core_keymem_U1143 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[711]), .Y(aes_core_keymem_n1515) );
  OAI2BB2X1 aes_core_keymem_U1142 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[710]), .Y(aes_core_keymem_n1527) );
  OAI2BB2X1 aes_core_keymem_U1141 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[709]), .Y(aes_core_keymem_n1539) );
  OAI2BB2X1 aes_core_keymem_U1140 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[708]), .Y(aes_core_keymem_n1551) );
  OAI2BB2X1 aes_core_keymem_U1139 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[707]), .Y(aes_core_keymem_n1563) );
  OAI2BB2X1 aes_core_keymem_U1138 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[706]), .Y(aes_core_keymem_n1575) );
  OAI2BB2X1 aes_core_keymem_U1137 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[705]), .Y(aes_core_keymem_n1587) );
  OAI2BB2X1 aes_core_keymem_U1136 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[704]), .Y(aes_core_keymem_n1599) );
  OAI2BB2X1 aes_core_keymem_U1135 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[703]), .Y(aes_core_keymem_n1611) );
  OAI2BB2X1 aes_core_keymem_U1134 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[702]), .Y(aes_core_keymem_n1623) );
  OAI2BB2X1 aes_core_keymem_U1133 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[701]), .Y(aes_core_keymem_n1635) );
  OAI2BB2X1 aes_core_keymem_U1132 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[700]), .Y(aes_core_keymem_n1647) );
  OAI2BB2X1 aes_core_keymem_U1131 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[699]), .Y(aes_core_keymem_n1659) );
  OAI2BB2X1 aes_core_keymem_U1130 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[698]), .Y(aes_core_keymem_n1671) );
  OAI2BB2X1 aes_core_keymem_U1129 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[697]), .Y(aes_core_keymem_n1683) );
  OAI2BB2X1 aes_core_keymem_U1128 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[696]), .Y(aes_core_keymem_n1695) );
  OAI2BB2X1 aes_core_keymem_U1127 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[695]), .Y(aes_core_keymem_n1707) );
  OAI2BB2X1 aes_core_keymem_U1126 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[694]), .Y(aes_core_keymem_n1719) );
  OAI2BB2X1 aes_core_keymem_U1125 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[693]), .Y(aes_core_keymem_n1731) );
  OAI2BB2X1 aes_core_keymem_U1124 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[692]), .Y(aes_core_keymem_n1743) );
  OAI2BB2X1 aes_core_keymem_U1123 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[691]), .Y(aes_core_keymem_n1755) );
  OAI2BB2X1 aes_core_keymem_U1122 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[690]), .Y(aes_core_keymem_n1767) );
  OAI2BB2X1 aes_core_keymem_U1121 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[689]), .Y(aes_core_keymem_n1779) );
  OAI2BB2X1 aes_core_keymem_U1120 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[688]), .Y(aes_core_keymem_n1791) );
  OAI2BB2X1 aes_core_keymem_U1119 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[687]), .Y(aes_core_keymem_n1803) );
  OAI2BB2X1 aes_core_keymem_U1118 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[686]), .Y(aes_core_keymem_n1815) );
  OAI2BB2X1 aes_core_keymem_U1117 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[685]), .Y(aes_core_keymem_n1827) );
  OAI2BB2X1 aes_core_keymem_U1116 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[684]), .Y(aes_core_keymem_n1839) );
  OAI2BB2X1 aes_core_keymem_U1115 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[683]), .Y(aes_core_keymem_n1851) );
  OAI2BB2X1 aes_core_keymem_U1114 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[682]), .Y(aes_core_keymem_n1863) );
  OAI2BB2X1 aes_core_keymem_U1113 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[681]), .Y(aes_core_keymem_n1875) );
  OAI2BB2X1 aes_core_keymem_U1112 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[680]), .Y(aes_core_keymem_n1887) );
  OAI2BB2X1 aes_core_keymem_U1111 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[679]), .Y(aes_core_keymem_n1899) );
  OAI2BB2X1 aes_core_keymem_U1110 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[678]), .Y(aes_core_keymem_n1911) );
  OAI2BB2X1 aes_core_keymem_U1109 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[677]), .Y(aes_core_keymem_n1923) );
  OAI2BB2X1 aes_core_keymem_U1108 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[676]), .Y(aes_core_keymem_n1935) );
  OAI2BB2X1 aes_core_keymem_U1107 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[675]), .Y(aes_core_keymem_n1947) );
  OAI2BB2X1 aes_core_keymem_U1106 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[674]), .Y(aes_core_keymem_n1959) );
  OAI2BB2X1 aes_core_keymem_U1105 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[673]), .Y(aes_core_keymem_n1971) );
  OAI2BB2X1 aes_core_keymem_U1104 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[672]), .Y(aes_core_keymem_n1983) );
  OAI2BB2X1 aes_core_keymem_U1103 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[671]), .Y(aes_core_keymem_n1995) );
  OAI2BB2X1 aes_core_keymem_U1102 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[670]), .Y(aes_core_keymem_n2007) );
  OAI2BB2X1 aes_core_keymem_U1101 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[669]), .Y(aes_core_keymem_n2019) );
  OAI2BB2X1 aes_core_keymem_U1100 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[668]), .Y(aes_core_keymem_n2031) );
  OAI2BB2X1 aes_core_keymem_U1099 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[667]), .Y(aes_core_keymem_n2043) );
  OAI2BB2X1 aes_core_keymem_U1098 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[666]), .Y(aes_core_keymem_n2055) );
  OAI2BB2X1 aes_core_keymem_U1097 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[665]), .Y(aes_core_keymem_n2067) );
  OAI2BB2X1 aes_core_keymem_U1096 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[664]), .Y(aes_core_keymem_n2079) );
  OAI2BB2X1 aes_core_keymem_U1095 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[663]), .Y(aes_core_keymem_n2091) );
  OAI2BB2X1 aes_core_keymem_U1094 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[662]), .Y(aes_core_keymem_n2103) );
  OAI2BB2X1 aes_core_keymem_U1093 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[661]), .Y(aes_core_keymem_n2115) );
  OAI2BB2X1 aes_core_keymem_U1092 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[660]), .Y(aes_core_keymem_n2127) );
  OAI2BB2X1 aes_core_keymem_U1091 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[659]), .Y(aes_core_keymem_n2139) );
  OAI2BB2X1 aes_core_keymem_U1090 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[658]), .Y(aes_core_keymem_n2151) );
  OAI2BB2X1 aes_core_keymem_U1089 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[657]), .Y(aes_core_keymem_n2163) );
  OAI2BB2X1 aes_core_keymem_U1088 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[656]), .Y(aes_core_keymem_n2175) );
  OAI2BB2X1 aes_core_keymem_U1087 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[655]), .Y(aes_core_keymem_n2187) );
  OAI2BB2X1 aes_core_keymem_U1086 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[654]), .Y(aes_core_keymem_n2199) );
  OAI2BB2X1 aes_core_keymem_U1085 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[653]), .Y(aes_core_keymem_n2211) );
  OAI2BB2X1 aes_core_keymem_U1084 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[652]), .Y(aes_core_keymem_n2223) );
  OAI2BB2X1 aes_core_keymem_U1083 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[651]), .Y(aes_core_keymem_n2235) );
  OAI2BB2X1 aes_core_keymem_U1082 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[650]), .Y(aes_core_keymem_n2247) );
  OAI2BB2X1 aes_core_keymem_U1081 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[649]), .Y(aes_core_keymem_n2259) );
  OAI2BB2X1 aes_core_keymem_U1080 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[648]), .Y(aes_core_keymem_n2271) );
  OAI2BB2X1 aes_core_keymem_U1079 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[647]), .Y(aes_core_keymem_n2283) );
  OAI2BB2X1 aes_core_keymem_U1078 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[646]), .Y(aes_core_keymem_n2295) );
  OAI2BB2X1 aes_core_keymem_U1077 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[645]), .Y(aes_core_keymem_n2307) );
  OAI2BB2X1 aes_core_keymem_U1076 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[644]), .Y(aes_core_keymem_n2319) );
  OAI2BB2X1 aes_core_keymem_U1075 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[643]), .Y(aes_core_keymem_n2331) );
  OAI2BB2X1 aes_core_keymem_U1074 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[642]), .Y(aes_core_keymem_n2343) );
  OAI2BB2X1 aes_core_keymem_U1073 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[641]), .Y(aes_core_keymem_n2355) );
  OAI2BB2X1 aes_core_keymem_U1072 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n548), .A0N(aes_core_keymem_n548), .A1N(
        aes_core_keymem_key_mem[640]), .Y(aes_core_keymem_n2367) );
  OAI2BB2X1 aes_core_keymem_U1071 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[255]), .Y(aes_core_keymem_n846) );
  OAI2BB2X1 aes_core_keymem_U1070 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[254]), .Y(aes_core_keymem_n858) );
  OAI2BB2X1 aes_core_keymem_U1069 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[253]), .Y(aes_core_keymem_n870) );
  OAI2BB2X1 aes_core_keymem_U1068 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[252]), .Y(aes_core_keymem_n882) );
  OAI2BB2X1 aes_core_keymem_U1067 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[251]), .Y(aes_core_keymem_n894) );
  OAI2BB2X1 aes_core_keymem_U1066 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[250]), .Y(aes_core_keymem_n906) );
  OAI2BB2X1 aes_core_keymem_U1065 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[249]), .Y(aes_core_keymem_n918) );
  OAI2BB2X1 aes_core_keymem_U1064 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[248]), .Y(aes_core_keymem_n930) );
  OAI2BB2X1 aes_core_keymem_U1063 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[247]), .Y(aes_core_keymem_n942) );
  OAI2BB2X1 aes_core_keymem_U1062 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[246]), .Y(aes_core_keymem_n954) );
  OAI2BB2X1 aes_core_keymem_U1061 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[245]), .Y(aes_core_keymem_n966) );
  OAI2BB2X1 aes_core_keymem_U1060 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[244]), .Y(aes_core_keymem_n978) );
  OAI2BB2X1 aes_core_keymem_U1059 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[243]), .Y(aes_core_keymem_n990) );
  OAI2BB2X1 aes_core_keymem_U1058 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[242]), .Y(aes_core_keymem_n1002) );
  OAI2BB2X1 aes_core_keymem_U1057 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[241]), .Y(aes_core_keymem_n1014) );
  OAI2BB2X1 aes_core_keymem_U1056 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[240]), .Y(aes_core_keymem_n1026) );
  OAI2BB2X1 aes_core_keymem_U1055 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[239]), .Y(aes_core_keymem_n1038) );
  OAI2BB2X1 aes_core_keymem_U1054 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[238]), .Y(aes_core_keymem_n1050) );
  OAI2BB2X1 aes_core_keymem_U1053 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[237]), .Y(aes_core_keymem_n1062) );
  OAI2BB2X1 aes_core_keymem_U1052 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[236]), .Y(aes_core_keymem_n1074) );
  OAI2BB2X1 aes_core_keymem_U1051 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[235]), .Y(aes_core_keymem_n1086) );
  OAI2BB2X1 aes_core_keymem_U1050 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[234]), .Y(aes_core_keymem_n1098) );
  OAI2BB2X1 aes_core_keymem_U1049 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[233]), .Y(aes_core_keymem_n1110) );
  OAI2BB2X1 aes_core_keymem_U1048 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[232]), .Y(aes_core_keymem_n1122) );
  OAI2BB2X1 aes_core_keymem_U1047 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[231]), .Y(aes_core_keymem_n1134) );
  OAI2BB2X1 aes_core_keymem_U1046 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[230]), .Y(aes_core_keymem_n1146) );
  OAI2BB2X1 aes_core_keymem_U1045 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[229]), .Y(aes_core_keymem_n1158) );
  OAI2BB2X1 aes_core_keymem_U1044 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[228]), .Y(aes_core_keymem_n1170) );
  OAI2BB2X1 aes_core_keymem_U1043 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[227]), .Y(aes_core_keymem_n1182) );
  OAI2BB2X1 aes_core_keymem_U1042 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[226]), .Y(aes_core_keymem_n1194) );
  OAI2BB2X1 aes_core_keymem_U1041 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[225]), .Y(aes_core_keymem_n1206) );
  OAI2BB2X1 aes_core_keymem_U1040 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[224]), .Y(aes_core_keymem_n1218) );
  OAI2BB2X1 aes_core_keymem_U1039 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[223]), .Y(aes_core_keymem_n1230) );
  OAI2BB2X1 aes_core_keymem_U1038 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[222]), .Y(aes_core_keymem_n1242) );
  OAI2BB2X1 aes_core_keymem_U1037 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[221]), .Y(aes_core_keymem_n1254) );
  OAI2BB2X1 aes_core_keymem_U1036 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[220]), .Y(aes_core_keymem_n1266) );
  OAI2BB2X1 aes_core_keymem_U1035 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[219]), .Y(aes_core_keymem_n1278) );
  OAI2BB2X1 aes_core_keymem_U1034 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[218]), .Y(aes_core_keymem_n1290) );
  OAI2BB2X1 aes_core_keymem_U1033 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[217]), .Y(aes_core_keymem_n1302) );
  OAI2BB2X1 aes_core_keymem_U1032 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[216]), .Y(aes_core_keymem_n1314) );
  OAI2BB2X1 aes_core_keymem_U1031 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[215]), .Y(aes_core_keymem_n1326) );
  OAI2BB2X1 aes_core_keymem_U1030 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[214]), .Y(aes_core_keymem_n1338) );
  OAI2BB2X1 aes_core_keymem_U1029 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[213]), .Y(aes_core_keymem_n1350) );
  OAI2BB2X1 aes_core_keymem_U1028 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[212]), .Y(aes_core_keymem_n1362) );
  OAI2BB2X1 aes_core_keymem_U1027 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[211]), .Y(aes_core_keymem_n1374) );
  OAI2BB2X1 aes_core_keymem_U1026 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[210]), .Y(aes_core_keymem_n1386) );
  OAI2BB2X1 aes_core_keymem_U1025 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[209]), .Y(aes_core_keymem_n1398) );
  OAI2BB2X1 aes_core_keymem_U1024 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[208]), .Y(aes_core_keymem_n1410) );
  OAI2BB2X1 aes_core_keymem_U1023 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[207]), .Y(aes_core_keymem_n1422) );
  OAI2BB2X1 aes_core_keymem_U1022 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[206]), .Y(aes_core_keymem_n1434) );
  OAI2BB2X1 aes_core_keymem_U1021 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[205]), .Y(aes_core_keymem_n1446) );
  OAI2BB2X1 aes_core_keymem_U1020 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[204]), .Y(aes_core_keymem_n1458) );
  OAI2BB2X1 aes_core_keymem_U1019 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[203]), .Y(aes_core_keymem_n1470) );
  OAI2BB2X1 aes_core_keymem_U1018 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[202]), .Y(aes_core_keymem_n1482) );
  OAI2BB2X1 aes_core_keymem_U1017 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[201]), .Y(aes_core_keymem_n1494) );
  OAI2BB2X1 aes_core_keymem_U1016 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[200]), .Y(aes_core_keymem_n1506) );
  OAI2BB2X1 aes_core_keymem_U1015 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[199]), .Y(aes_core_keymem_n1518) );
  OAI2BB2X1 aes_core_keymem_U1014 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[198]), .Y(aes_core_keymem_n1530) );
  OAI2BB2X1 aes_core_keymem_U1013 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[197]), .Y(aes_core_keymem_n1542) );
  OAI2BB2X1 aes_core_keymem_U1012 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[196]), .Y(aes_core_keymem_n1554) );
  OAI2BB2X1 aes_core_keymem_U1011 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[195]), .Y(aes_core_keymem_n1566) );
  OAI2BB2X1 aes_core_keymem_U1010 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[194]), .Y(aes_core_keymem_n1578) );
  OAI2BB2X1 aes_core_keymem_U1009 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[193]), .Y(aes_core_keymem_n1590) );
  OAI2BB2X1 aes_core_keymem_U1008 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[192]), .Y(aes_core_keymem_n1602) );
  OAI2BB2X1 aes_core_keymem_U1007 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[191]), .Y(aes_core_keymem_n1614) );
  OAI2BB2X1 aes_core_keymem_U1006 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[190]), .Y(aes_core_keymem_n1626) );
  OAI2BB2X1 aes_core_keymem_U1005 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[189]), .Y(aes_core_keymem_n1638) );
  OAI2BB2X1 aes_core_keymem_U1004 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[188]), .Y(aes_core_keymem_n1650) );
  OAI2BB2X1 aes_core_keymem_U1003 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[187]), .Y(aes_core_keymem_n1662) );
  OAI2BB2X1 aes_core_keymem_U1002 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[186]), .Y(aes_core_keymem_n1674) );
  OAI2BB2X1 aes_core_keymem_U1001 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[185]), .Y(aes_core_keymem_n1686) );
  OAI2BB2X1 aes_core_keymem_U1000 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[184]), .Y(aes_core_keymem_n1698) );
  OAI2BB2X1 aes_core_keymem_U999 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[183]), .Y(aes_core_keymem_n1710) );
  OAI2BB2X1 aes_core_keymem_U998 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[182]), .Y(aes_core_keymem_n1722) );
  OAI2BB2X1 aes_core_keymem_U997 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[181]), .Y(aes_core_keymem_n1734) );
  OAI2BB2X1 aes_core_keymem_U996 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[180]), .Y(aes_core_keymem_n1746) );
  OAI2BB2X1 aes_core_keymem_U995 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[179]), .Y(aes_core_keymem_n1758) );
  OAI2BB2X1 aes_core_keymem_U994 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[178]), .Y(aes_core_keymem_n1770) );
  OAI2BB2X1 aes_core_keymem_U993 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[177]), .Y(aes_core_keymem_n1782) );
  OAI2BB2X1 aes_core_keymem_U992 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[176]), .Y(aes_core_keymem_n1794) );
  OAI2BB2X1 aes_core_keymem_U991 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[175]), .Y(aes_core_keymem_n1806) );
  OAI2BB2X1 aes_core_keymem_U990 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[174]), .Y(aes_core_keymem_n1818) );
  OAI2BB2X1 aes_core_keymem_U989 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[173]), .Y(aes_core_keymem_n1830) );
  OAI2BB2X1 aes_core_keymem_U988 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[172]), .Y(aes_core_keymem_n1842) );
  OAI2BB2X1 aes_core_keymem_U987 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[171]), .Y(aes_core_keymem_n1854) );
  OAI2BB2X1 aes_core_keymem_U986 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[170]), .Y(aes_core_keymem_n1866) );
  OAI2BB2X1 aes_core_keymem_U985 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[169]), .Y(aes_core_keymem_n1878) );
  OAI2BB2X1 aes_core_keymem_U984 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[168]), .Y(aes_core_keymem_n1890) );
  OAI2BB2X1 aes_core_keymem_U983 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[167]), .Y(aes_core_keymem_n1902) );
  OAI2BB2X1 aes_core_keymem_U982 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[166]), .Y(aes_core_keymem_n1914) );
  OAI2BB2X1 aes_core_keymem_U981 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[165]), .Y(aes_core_keymem_n1926) );
  OAI2BB2X1 aes_core_keymem_U980 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[164]), .Y(aes_core_keymem_n1938) );
  OAI2BB2X1 aes_core_keymem_U979 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[163]), .Y(aes_core_keymem_n1950) );
  OAI2BB2X1 aes_core_keymem_U978 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[162]), .Y(aes_core_keymem_n1962) );
  OAI2BB2X1 aes_core_keymem_U977 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[161]), .Y(aes_core_keymem_n1974) );
  OAI2BB2X1 aes_core_keymem_U976 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[160]), .Y(aes_core_keymem_n1986) );
  OAI2BB2X1 aes_core_keymem_U975 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[159]), .Y(aes_core_keymem_n1998) );
  OAI2BB2X1 aes_core_keymem_U974 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[158]), .Y(aes_core_keymem_n2010) );
  OAI2BB2X1 aes_core_keymem_U973 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[157]), .Y(aes_core_keymem_n2022) );
  OAI2BB2X1 aes_core_keymem_U972 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[156]), .Y(aes_core_keymem_n2034) );
  OAI2BB2X1 aes_core_keymem_U971 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[155]), .Y(aes_core_keymem_n2046) );
  OAI2BB2X1 aes_core_keymem_U970 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[154]), .Y(aes_core_keymem_n2058) );
  OAI2BB2X1 aes_core_keymem_U969 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[153]), .Y(aes_core_keymem_n2070) );
  OAI2BB2X1 aes_core_keymem_U968 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[152]), .Y(aes_core_keymem_n2082) );
  OAI2BB2X1 aes_core_keymem_U967 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[151]), .Y(aes_core_keymem_n2094) );
  OAI2BB2X1 aes_core_keymem_U966 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[150]), .Y(aes_core_keymem_n2106) );
  OAI2BB2X1 aes_core_keymem_U965 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[149]), .Y(aes_core_keymem_n2118) );
  OAI2BB2X1 aes_core_keymem_U964 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[148]), .Y(aes_core_keymem_n2130) );
  OAI2BB2X1 aes_core_keymem_U963 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[147]), .Y(aes_core_keymem_n2142) );
  OAI2BB2X1 aes_core_keymem_U962 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[146]), .Y(aes_core_keymem_n2154) );
  OAI2BB2X1 aes_core_keymem_U961 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[145]), .Y(aes_core_keymem_n2166) );
  OAI2BB2X1 aes_core_keymem_U960 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[144]), .Y(aes_core_keymem_n2178) );
  OAI2BB2X1 aes_core_keymem_U959 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[143]), .Y(aes_core_keymem_n2190) );
  OAI2BB2X1 aes_core_keymem_U958 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[142]), .Y(aes_core_keymem_n2202) );
  OAI2BB2X1 aes_core_keymem_U957 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[141]), .Y(aes_core_keymem_n2214) );
  OAI2BB2X1 aes_core_keymem_U956 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[140]), .Y(aes_core_keymem_n2226) );
  OAI2BB2X1 aes_core_keymem_U955 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[139]), .Y(aes_core_keymem_n2238) );
  OAI2BB2X1 aes_core_keymem_U954 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[138]), .Y(aes_core_keymem_n2250) );
  OAI2BB2X1 aes_core_keymem_U953 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[137]), .Y(aes_core_keymem_n2262) );
  OAI2BB2X1 aes_core_keymem_U952 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[136]), .Y(aes_core_keymem_n2274) );
  OAI2BB2X1 aes_core_keymem_U951 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[135]), .Y(aes_core_keymem_n2286) );
  OAI2BB2X1 aes_core_keymem_U950 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[134]), .Y(aes_core_keymem_n2298) );
  OAI2BB2X1 aes_core_keymem_U949 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[133]), .Y(aes_core_keymem_n2310) );
  OAI2BB2X1 aes_core_keymem_U948 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[132]), .Y(aes_core_keymem_n2322) );
  OAI2BB2X1 aes_core_keymem_U947 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[131]), .Y(aes_core_keymem_n2334) );
  OAI2BB2X1 aes_core_keymem_U946 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[130]), .Y(aes_core_keymem_n2346) );
  OAI2BB2X1 aes_core_keymem_U945 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[129]), .Y(aes_core_keymem_n2358) );
  OAI2BB2X1 aes_core_keymem_U944 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n551), .A0N(aes_core_keymem_n551), .A1N(
        aes_core_keymem_key_mem[128]), .Y(aes_core_keymem_n2370) );
  OAI2BB2X1 aes_core_keymem_U943 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[511]), .Y(aes_core_keymem_n848) );
  OAI2BB2X1 aes_core_keymem_U942 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[510]), .Y(aes_core_keymem_n860) );
  OAI2BB2X1 aes_core_keymem_U941 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[509]), .Y(aes_core_keymem_n872) );
  OAI2BB2X1 aes_core_keymem_U940 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[508]), .Y(aes_core_keymem_n884) );
  OAI2BB2X1 aes_core_keymem_U939 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[507]), .Y(aes_core_keymem_n896) );
  OAI2BB2X1 aes_core_keymem_U938 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[506]), .Y(aes_core_keymem_n908) );
  OAI2BB2X1 aes_core_keymem_U937 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[505]), .Y(aes_core_keymem_n920) );
  OAI2BB2X1 aes_core_keymem_U936 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[504]), .Y(aes_core_keymem_n932) );
  OAI2BB2X1 aes_core_keymem_U935 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[503]), .Y(aes_core_keymem_n944) );
  OAI2BB2X1 aes_core_keymem_U934 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[502]), .Y(aes_core_keymem_n956) );
  OAI2BB2X1 aes_core_keymem_U933 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[501]), .Y(aes_core_keymem_n968) );
  OAI2BB2X1 aes_core_keymem_U932 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[500]), .Y(aes_core_keymem_n980) );
  OAI2BB2X1 aes_core_keymem_U931 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[499]), .Y(aes_core_keymem_n992) );
  OAI2BB2X1 aes_core_keymem_U930 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[498]), .Y(aes_core_keymem_n1004) );
  OAI2BB2X1 aes_core_keymem_U929 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[497]), .Y(aes_core_keymem_n1016) );
  OAI2BB2X1 aes_core_keymem_U928 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[496]), .Y(aes_core_keymem_n1028) );
  OAI2BB2X1 aes_core_keymem_U927 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[495]), .Y(aes_core_keymem_n1040) );
  OAI2BB2X1 aes_core_keymem_U926 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[494]), .Y(aes_core_keymem_n1052) );
  OAI2BB2X1 aes_core_keymem_U925 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[493]), .Y(aes_core_keymem_n1064) );
  OAI2BB2X1 aes_core_keymem_U924 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[492]), .Y(aes_core_keymem_n1076) );
  OAI2BB2X1 aes_core_keymem_U923 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[491]), .Y(aes_core_keymem_n1088) );
  OAI2BB2X1 aes_core_keymem_U922 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[490]), .Y(aes_core_keymem_n1100) );
  OAI2BB2X1 aes_core_keymem_U921 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[489]), .Y(aes_core_keymem_n1112) );
  OAI2BB2X1 aes_core_keymem_U920 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[488]), .Y(aes_core_keymem_n1124) );
  OAI2BB2X1 aes_core_keymem_U919 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[487]), .Y(aes_core_keymem_n1136) );
  OAI2BB2X1 aes_core_keymem_U918 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[486]), .Y(aes_core_keymem_n1148) );
  OAI2BB2X1 aes_core_keymem_U917 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[485]), .Y(aes_core_keymem_n1160) );
  OAI2BB2X1 aes_core_keymem_U916 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[484]), .Y(aes_core_keymem_n1172) );
  OAI2BB2X1 aes_core_keymem_U915 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[483]), .Y(aes_core_keymem_n1184) );
  OAI2BB2X1 aes_core_keymem_U914 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[482]), .Y(aes_core_keymem_n1196) );
  OAI2BB2X1 aes_core_keymem_U913 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[481]), .Y(aes_core_keymem_n1208) );
  OAI2BB2X1 aes_core_keymem_U912 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[480]), .Y(aes_core_keymem_n1220) );
  OAI2BB2X1 aes_core_keymem_U911 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[479]), .Y(aes_core_keymem_n1232) );
  OAI2BB2X1 aes_core_keymem_U910 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[478]), .Y(aes_core_keymem_n1244) );
  OAI2BB2X1 aes_core_keymem_U909 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[477]), .Y(aes_core_keymem_n1256) );
  OAI2BB2X1 aes_core_keymem_U908 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[476]), .Y(aes_core_keymem_n1268) );
  OAI2BB2X1 aes_core_keymem_U907 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[475]), .Y(aes_core_keymem_n1280) );
  OAI2BB2X1 aes_core_keymem_U906 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[474]), .Y(aes_core_keymem_n1292) );
  OAI2BB2X1 aes_core_keymem_U905 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[473]), .Y(aes_core_keymem_n1304) );
  OAI2BB2X1 aes_core_keymem_U904 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[472]), .Y(aes_core_keymem_n1316) );
  OAI2BB2X1 aes_core_keymem_U903 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[471]), .Y(aes_core_keymem_n1328) );
  OAI2BB2X1 aes_core_keymem_U902 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[470]), .Y(aes_core_keymem_n1340) );
  OAI2BB2X1 aes_core_keymem_U901 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[469]), .Y(aes_core_keymem_n1352) );
  OAI2BB2X1 aes_core_keymem_U900 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[468]), .Y(aes_core_keymem_n1364) );
  OAI2BB2X1 aes_core_keymem_U899 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[467]), .Y(aes_core_keymem_n1376) );
  OAI2BB2X1 aes_core_keymem_U898 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[466]), .Y(aes_core_keymem_n1388) );
  OAI2BB2X1 aes_core_keymem_U897 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[465]), .Y(aes_core_keymem_n1400) );
  OAI2BB2X1 aes_core_keymem_U896 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[464]), .Y(aes_core_keymem_n1412) );
  OAI2BB2X1 aes_core_keymem_U895 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[463]), .Y(aes_core_keymem_n1424) );
  OAI2BB2X1 aes_core_keymem_U894 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[462]), .Y(aes_core_keymem_n1436) );
  OAI2BB2X1 aes_core_keymem_U893 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[461]), .Y(aes_core_keymem_n1448) );
  OAI2BB2X1 aes_core_keymem_U892 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[460]), .Y(aes_core_keymem_n1460) );
  OAI2BB2X1 aes_core_keymem_U891 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[459]), .Y(aes_core_keymem_n1472) );
  OAI2BB2X1 aes_core_keymem_U890 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[458]), .Y(aes_core_keymem_n1484) );
  OAI2BB2X1 aes_core_keymem_U889 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[457]), .Y(aes_core_keymem_n1496) );
  OAI2BB2X1 aes_core_keymem_U888 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[456]), .Y(aes_core_keymem_n1508) );
  OAI2BB2X1 aes_core_keymem_U887 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[455]), .Y(aes_core_keymem_n1520) );
  OAI2BB2X1 aes_core_keymem_U886 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[454]), .Y(aes_core_keymem_n1532) );
  OAI2BB2X1 aes_core_keymem_U885 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[453]), .Y(aes_core_keymem_n1544) );
  OAI2BB2X1 aes_core_keymem_U884 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[452]), .Y(aes_core_keymem_n1556) );
  OAI2BB2X1 aes_core_keymem_U883 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[451]), .Y(aes_core_keymem_n1568) );
  OAI2BB2X1 aes_core_keymem_U882 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[450]), .Y(aes_core_keymem_n1580) );
  OAI2BB2X1 aes_core_keymem_U881 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[449]), .Y(aes_core_keymem_n1592) );
  OAI2BB2X1 aes_core_keymem_U880 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[448]), .Y(aes_core_keymem_n1604) );
  OAI2BB2X1 aes_core_keymem_U879 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[447]), .Y(aes_core_keymem_n1616) );
  OAI2BB2X1 aes_core_keymem_U878 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[446]), .Y(aes_core_keymem_n1628) );
  OAI2BB2X1 aes_core_keymem_U877 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[445]), .Y(aes_core_keymem_n1640) );
  OAI2BB2X1 aes_core_keymem_U876 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[444]), .Y(aes_core_keymem_n1652) );
  OAI2BB2X1 aes_core_keymem_U875 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[443]), .Y(aes_core_keymem_n1664) );
  OAI2BB2X1 aes_core_keymem_U874 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[442]), .Y(aes_core_keymem_n1676) );
  OAI2BB2X1 aes_core_keymem_U873 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[441]), .Y(aes_core_keymem_n1688) );
  OAI2BB2X1 aes_core_keymem_U872 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[440]), .Y(aes_core_keymem_n1700) );
  OAI2BB2X1 aes_core_keymem_U871 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[439]), .Y(aes_core_keymem_n1712) );
  OAI2BB2X1 aes_core_keymem_U870 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[438]), .Y(aes_core_keymem_n1724) );
  OAI2BB2X1 aes_core_keymem_U869 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[437]), .Y(aes_core_keymem_n1736) );
  OAI2BB2X1 aes_core_keymem_U868 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[436]), .Y(aes_core_keymem_n1748) );
  OAI2BB2X1 aes_core_keymem_U867 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[435]), .Y(aes_core_keymem_n1760) );
  OAI2BB2X1 aes_core_keymem_U866 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[434]), .Y(aes_core_keymem_n1772) );
  OAI2BB2X1 aes_core_keymem_U865 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[433]), .Y(aes_core_keymem_n1784) );
  OAI2BB2X1 aes_core_keymem_U864 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[432]), .Y(aes_core_keymem_n1796) );
  OAI2BB2X1 aes_core_keymem_U863 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[431]), .Y(aes_core_keymem_n1808) );
  OAI2BB2X1 aes_core_keymem_U862 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[430]), .Y(aes_core_keymem_n1820) );
  OAI2BB2X1 aes_core_keymem_U861 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[429]), .Y(aes_core_keymem_n1832) );
  OAI2BB2X1 aes_core_keymem_U860 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[428]), .Y(aes_core_keymem_n1844) );
  OAI2BB2X1 aes_core_keymem_U859 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[427]), .Y(aes_core_keymem_n1856) );
  OAI2BB2X1 aes_core_keymem_U858 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[426]), .Y(aes_core_keymem_n1868) );
  OAI2BB2X1 aes_core_keymem_U857 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[425]), .Y(aes_core_keymem_n1880) );
  OAI2BB2X1 aes_core_keymem_U856 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[424]), .Y(aes_core_keymem_n1892) );
  OAI2BB2X1 aes_core_keymem_U855 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[423]), .Y(aes_core_keymem_n1904) );
  OAI2BB2X1 aes_core_keymem_U854 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[422]), .Y(aes_core_keymem_n1916) );
  OAI2BB2X1 aes_core_keymem_U853 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[421]), .Y(aes_core_keymem_n1928) );
  OAI2BB2X1 aes_core_keymem_U852 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[420]), .Y(aes_core_keymem_n1940) );
  OAI2BB2X1 aes_core_keymem_U851 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[419]), .Y(aes_core_keymem_n1952) );
  OAI2BB2X1 aes_core_keymem_U850 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[418]), .Y(aes_core_keymem_n1964) );
  OAI2BB2X1 aes_core_keymem_U849 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[417]), .Y(aes_core_keymem_n1976) );
  OAI2BB2X1 aes_core_keymem_U848 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[416]), .Y(aes_core_keymem_n1988) );
  OAI2BB2X1 aes_core_keymem_U847 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[415]), .Y(aes_core_keymem_n2000) );
  OAI2BB2X1 aes_core_keymem_U846 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[414]), .Y(aes_core_keymem_n2012) );
  OAI2BB2X1 aes_core_keymem_U845 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[413]), .Y(aes_core_keymem_n2024) );
  OAI2BB2X1 aes_core_keymem_U844 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[412]), .Y(aes_core_keymem_n2036) );
  OAI2BB2X1 aes_core_keymem_U843 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[411]), .Y(aes_core_keymem_n2048) );
  OAI2BB2X1 aes_core_keymem_U842 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[410]), .Y(aes_core_keymem_n2060) );
  OAI2BB2X1 aes_core_keymem_U841 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[409]), .Y(aes_core_keymem_n2072) );
  OAI2BB2X1 aes_core_keymem_U840 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[408]), .Y(aes_core_keymem_n2084) );
  OAI2BB2X1 aes_core_keymem_U839 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[407]), .Y(aes_core_keymem_n2096) );
  OAI2BB2X1 aes_core_keymem_U838 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[406]), .Y(aes_core_keymem_n2108) );
  OAI2BB2X1 aes_core_keymem_U837 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[405]), .Y(aes_core_keymem_n2120) );
  OAI2BB2X1 aes_core_keymem_U836 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[404]), .Y(aes_core_keymem_n2132) );
  OAI2BB2X1 aes_core_keymem_U835 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[403]), .Y(aes_core_keymem_n2144) );
  OAI2BB2X1 aes_core_keymem_U834 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[402]), .Y(aes_core_keymem_n2156) );
  OAI2BB2X1 aes_core_keymem_U833 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[401]), .Y(aes_core_keymem_n2168) );
  OAI2BB2X1 aes_core_keymem_U832 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[400]), .Y(aes_core_keymem_n2180) );
  OAI2BB2X1 aes_core_keymem_U831 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[399]), .Y(aes_core_keymem_n2192) );
  OAI2BB2X1 aes_core_keymem_U830 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[398]), .Y(aes_core_keymem_n2204) );
  OAI2BB2X1 aes_core_keymem_U829 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[397]), .Y(aes_core_keymem_n2216) );
  OAI2BB2X1 aes_core_keymem_U828 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[396]), .Y(aes_core_keymem_n2228) );
  OAI2BB2X1 aes_core_keymem_U827 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[395]), .Y(aes_core_keymem_n2240) );
  OAI2BB2X1 aes_core_keymem_U826 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[394]), .Y(aes_core_keymem_n2252) );
  OAI2BB2X1 aes_core_keymem_U825 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[393]), .Y(aes_core_keymem_n2264) );
  OAI2BB2X1 aes_core_keymem_U824 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[392]), .Y(aes_core_keymem_n2276) );
  OAI2BB2X1 aes_core_keymem_U823 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[391]), .Y(aes_core_keymem_n2288) );
  OAI2BB2X1 aes_core_keymem_U822 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[390]), .Y(aes_core_keymem_n2300) );
  OAI2BB2X1 aes_core_keymem_U821 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[389]), .Y(aes_core_keymem_n2312) );
  OAI2BB2X1 aes_core_keymem_U820 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[388]), .Y(aes_core_keymem_n2324) );
  OAI2BB2X1 aes_core_keymem_U819 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[387]), .Y(aes_core_keymem_n2336) );
  OAI2BB2X1 aes_core_keymem_U818 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[386]), .Y(aes_core_keymem_n2348) );
  OAI2BB2X1 aes_core_keymem_U817 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[385]), .Y(aes_core_keymem_n2360) );
  OAI2BB2X1 aes_core_keymem_U816 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n553), .A0N(aes_core_keymem_n553), .A1N(
        aes_core_keymem_key_mem[384]), .Y(aes_core_keymem_n2372) );
  OAI2BB2X1 aes_core_keymem_U815 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[127]), .Y(aes_core_keymem_n845) );
  OAI2BB2X1 aes_core_keymem_U814 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[126]), .Y(aes_core_keymem_n857) );
  OAI2BB2X1 aes_core_keymem_U813 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[125]), .Y(aes_core_keymem_n869) );
  OAI2BB2X1 aes_core_keymem_U812 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[124]), .Y(aes_core_keymem_n881) );
  OAI2BB2X1 aes_core_keymem_U811 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[123]), .Y(aes_core_keymem_n893) );
  OAI2BB2X1 aes_core_keymem_U810 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[122]), .Y(aes_core_keymem_n905) );
  OAI2BB2X1 aes_core_keymem_U809 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[121]), .Y(aes_core_keymem_n917) );
  OAI2BB2X1 aes_core_keymem_U808 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[120]), .Y(aes_core_keymem_n929) );
  OAI2BB2X1 aes_core_keymem_U807 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[119]), .Y(aes_core_keymem_n941) );
  OAI2BB2X1 aes_core_keymem_U806 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[118]), .Y(aes_core_keymem_n953) );
  OAI2BB2X1 aes_core_keymem_U805 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[117]), .Y(aes_core_keymem_n965) );
  OAI2BB2X1 aes_core_keymem_U804 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[116]), .Y(aes_core_keymem_n977) );
  OAI2BB2X1 aes_core_keymem_U803 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[115]), .Y(aes_core_keymem_n989) );
  OAI2BB2X1 aes_core_keymem_U802 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[114]), .Y(aes_core_keymem_n1001) );
  OAI2BB2X1 aes_core_keymem_U801 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[113]), .Y(aes_core_keymem_n1013) );
  OAI2BB2X1 aes_core_keymem_U800 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[112]), .Y(aes_core_keymem_n1025) );
  OAI2BB2X1 aes_core_keymem_U799 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[111]), .Y(aes_core_keymem_n1037) );
  OAI2BB2X1 aes_core_keymem_U798 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[110]), .Y(aes_core_keymem_n1049) );
  OAI2BB2X1 aes_core_keymem_U797 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[109]), .Y(aes_core_keymem_n1061) );
  OAI2BB2X1 aes_core_keymem_U796 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[108]), .Y(aes_core_keymem_n1073) );
  OAI2BB2X1 aes_core_keymem_U795 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[107]), .Y(aes_core_keymem_n1085) );
  OAI2BB2X1 aes_core_keymem_U794 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[106]), .Y(aes_core_keymem_n1097) );
  OAI2BB2X1 aes_core_keymem_U793 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[105]), .Y(aes_core_keymem_n1109) );
  OAI2BB2X1 aes_core_keymem_U792 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[104]), .Y(aes_core_keymem_n1121) );
  OAI2BB2X1 aes_core_keymem_U791 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[103]), .Y(aes_core_keymem_n1133) );
  OAI2BB2X1 aes_core_keymem_U790 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[102]), .Y(aes_core_keymem_n1145) );
  OAI2BB2X1 aes_core_keymem_U789 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[101]), .Y(aes_core_keymem_n1157) );
  OAI2BB2X1 aes_core_keymem_U788 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[100]), .Y(aes_core_keymem_n1169) );
  OAI2BB2X1 aes_core_keymem_U787 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[99]), .Y(aes_core_keymem_n1181) );
  OAI2BB2X1 aes_core_keymem_U786 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[98]), .Y(aes_core_keymem_n1193) );
  OAI2BB2X1 aes_core_keymem_U785 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[97]), .Y(aes_core_keymem_n1205) );
  OAI2BB2X1 aes_core_keymem_U784 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[96]), .Y(aes_core_keymem_n1217) );
  OAI2BB2X1 aes_core_keymem_U783 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[95]), .Y(aes_core_keymem_n1229) );
  OAI2BB2X1 aes_core_keymem_U782 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[94]), .Y(aes_core_keymem_n1241) );
  OAI2BB2X1 aes_core_keymem_U781 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[93]), .Y(aes_core_keymem_n1253) );
  OAI2BB2X1 aes_core_keymem_U780 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[92]), .Y(aes_core_keymem_n1265) );
  OAI2BB2X1 aes_core_keymem_U779 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[91]), .Y(aes_core_keymem_n1277) );
  OAI2BB2X1 aes_core_keymem_U778 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[90]), .Y(aes_core_keymem_n1289) );
  OAI2BB2X1 aes_core_keymem_U777 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[89]), .Y(aes_core_keymem_n1301) );
  OAI2BB2X1 aes_core_keymem_U776 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[88]), .Y(aes_core_keymem_n1313) );
  OAI2BB2X1 aes_core_keymem_U775 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[87]), .Y(aes_core_keymem_n1325) );
  OAI2BB2X1 aes_core_keymem_U774 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[86]), .Y(aes_core_keymem_n1337) );
  OAI2BB2X1 aes_core_keymem_U773 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[85]), .Y(aes_core_keymem_n1349) );
  OAI2BB2X1 aes_core_keymem_U772 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[84]), .Y(aes_core_keymem_n1361) );
  OAI2BB2X1 aes_core_keymem_U771 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[83]), .Y(aes_core_keymem_n1373) );
  OAI2BB2X1 aes_core_keymem_U770 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[82]), .Y(aes_core_keymem_n1385) );
  OAI2BB2X1 aes_core_keymem_U769 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[81]), .Y(aes_core_keymem_n1397) );
  OAI2BB2X1 aes_core_keymem_U768 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[80]), .Y(aes_core_keymem_n1409) );
  OAI2BB2X1 aes_core_keymem_U767 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[79]), .Y(aes_core_keymem_n1421) );
  OAI2BB2X1 aes_core_keymem_U766 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[78]), .Y(aes_core_keymem_n1433) );
  OAI2BB2X1 aes_core_keymem_U765 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[77]), .Y(aes_core_keymem_n1445) );
  OAI2BB2X1 aes_core_keymem_U764 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[76]), .Y(aes_core_keymem_n1457) );
  OAI2BB2X1 aes_core_keymem_U763 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[75]), .Y(aes_core_keymem_n1469) );
  OAI2BB2X1 aes_core_keymem_U762 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[74]), .Y(aes_core_keymem_n1481) );
  OAI2BB2X1 aes_core_keymem_U761 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[73]), .Y(aes_core_keymem_n1493) );
  OAI2BB2X1 aes_core_keymem_U760 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[72]), .Y(aes_core_keymem_n1505) );
  OAI2BB2X1 aes_core_keymem_U759 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[71]), .Y(aes_core_keymem_n1517) );
  OAI2BB2X1 aes_core_keymem_U758 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[70]), .Y(aes_core_keymem_n1529) );
  OAI2BB2X1 aes_core_keymem_U757 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[69]), .Y(aes_core_keymem_n1541) );
  OAI2BB2X1 aes_core_keymem_U756 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[68]), .Y(aes_core_keymem_n1553) );
  OAI2BB2X1 aes_core_keymem_U755 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[67]), .Y(aes_core_keymem_n1565) );
  OAI2BB2X1 aes_core_keymem_U754 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[66]), .Y(aes_core_keymem_n1577) );
  OAI2BB2X1 aes_core_keymem_U753 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[65]), .Y(aes_core_keymem_n1589) );
  OAI2BB2X1 aes_core_keymem_U752 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[64]), .Y(aes_core_keymem_n1601) );
  OAI2BB2X1 aes_core_keymem_U751 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[63]), .Y(aes_core_keymem_n1613) );
  OAI2BB2X1 aes_core_keymem_U750 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[62]), .Y(aes_core_keymem_n1625) );
  OAI2BB2X1 aes_core_keymem_U749 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[61]), .Y(aes_core_keymem_n1637) );
  OAI2BB2X1 aes_core_keymem_U748 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[60]), .Y(aes_core_keymem_n1649) );
  OAI2BB2X1 aes_core_keymem_U747 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[59]), .Y(aes_core_keymem_n1661) );
  OAI2BB2X1 aes_core_keymem_U746 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[58]), .Y(aes_core_keymem_n1673) );
  OAI2BB2X1 aes_core_keymem_U745 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[57]), .Y(aes_core_keymem_n1685) );
  OAI2BB2X1 aes_core_keymem_U744 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[56]), .Y(aes_core_keymem_n1697) );
  OAI2BB2X1 aes_core_keymem_U743 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[55]), .Y(aes_core_keymem_n1709) );
  OAI2BB2X1 aes_core_keymem_U742 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[54]), .Y(aes_core_keymem_n1721) );
  OAI2BB2X1 aes_core_keymem_U741 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[53]), .Y(aes_core_keymem_n1733) );
  OAI2BB2X1 aes_core_keymem_U740 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[52]), .Y(aes_core_keymem_n1745) );
  OAI2BB2X1 aes_core_keymem_U739 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[51]), .Y(aes_core_keymem_n1757) );
  OAI2BB2X1 aes_core_keymem_U738 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[50]), .Y(aes_core_keymem_n1769) );
  OAI2BB2X1 aes_core_keymem_U737 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[49]), .Y(aes_core_keymem_n1781) );
  OAI2BB2X1 aes_core_keymem_U736 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[48]), .Y(aes_core_keymem_n1793) );
  OAI2BB2X1 aes_core_keymem_U735 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[47]), .Y(aes_core_keymem_n1805) );
  OAI2BB2X1 aes_core_keymem_U734 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[46]), .Y(aes_core_keymem_n1817) );
  OAI2BB2X1 aes_core_keymem_U733 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[45]), .Y(aes_core_keymem_n1829) );
  OAI2BB2X1 aes_core_keymem_U732 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[44]), .Y(aes_core_keymem_n1841) );
  OAI2BB2X1 aes_core_keymem_U731 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[43]), .Y(aes_core_keymem_n1853) );
  OAI2BB2X1 aes_core_keymem_U730 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[42]), .Y(aes_core_keymem_n1865) );
  OAI2BB2X1 aes_core_keymem_U729 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[41]), .Y(aes_core_keymem_n1877) );
  OAI2BB2X1 aes_core_keymem_U728 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[40]), .Y(aes_core_keymem_n1889) );
  OAI2BB2X1 aes_core_keymem_U727 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[39]), .Y(aes_core_keymem_n1901) );
  OAI2BB2X1 aes_core_keymem_U726 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[38]), .Y(aes_core_keymem_n1913) );
  OAI2BB2X1 aes_core_keymem_U725 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[37]), .Y(aes_core_keymem_n1925) );
  OAI2BB2X1 aes_core_keymem_U724 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[36]), .Y(aes_core_keymem_n1937) );
  OAI2BB2X1 aes_core_keymem_U723 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[35]), .Y(aes_core_keymem_n1949) );
  OAI2BB2X1 aes_core_keymem_U722 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[34]), .Y(aes_core_keymem_n1961) );
  OAI2BB2X1 aes_core_keymem_U721 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[33]), .Y(aes_core_keymem_n1973) );
  OAI2BB2X1 aes_core_keymem_U720 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[32]), .Y(aes_core_keymem_n1985) );
  OAI2BB2X1 aes_core_keymem_U719 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[31]), .Y(aes_core_keymem_n1997) );
  OAI2BB2X1 aes_core_keymem_U718 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[30]), .Y(aes_core_keymem_n2009) );
  OAI2BB2X1 aes_core_keymem_U717 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[29]), .Y(aes_core_keymem_n2021) );
  OAI2BB2X1 aes_core_keymem_U716 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[28]), .Y(aes_core_keymem_n2033) );
  OAI2BB2X1 aes_core_keymem_U715 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[27]), .Y(aes_core_keymem_n2045) );
  OAI2BB2X1 aes_core_keymem_U714 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[26]), .Y(aes_core_keymem_n2057) );
  OAI2BB2X1 aes_core_keymem_U713 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[25]), .Y(aes_core_keymem_n2069) );
  OAI2BB2X1 aes_core_keymem_U712 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[24]), .Y(aes_core_keymem_n2081) );
  OAI2BB2X1 aes_core_keymem_U711 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[23]), .Y(aes_core_keymem_n2093) );
  OAI2BB2X1 aes_core_keymem_U710 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[22]), .Y(aes_core_keymem_n2105) );
  OAI2BB2X1 aes_core_keymem_U709 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[21]), .Y(aes_core_keymem_n2117) );
  OAI2BB2X1 aes_core_keymem_U708 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[20]), .Y(aes_core_keymem_n2129) );
  OAI2BB2X1 aes_core_keymem_U707 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[19]), .Y(aes_core_keymem_n2141) );
  OAI2BB2X1 aes_core_keymem_U706 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[18]), .Y(aes_core_keymem_n2153) );
  OAI2BB2X1 aes_core_keymem_U705 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[17]), .Y(aes_core_keymem_n2165) );
  OAI2BB2X1 aes_core_keymem_U704 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[16]), .Y(aes_core_keymem_n2177) );
  OAI2BB2X1 aes_core_keymem_U703 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[15]), .Y(aes_core_keymem_n2189) );
  OAI2BB2X1 aes_core_keymem_U702 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[14]), .Y(aes_core_keymem_n2201) );
  OAI2BB2X1 aes_core_keymem_U701 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[13]), .Y(aes_core_keymem_n2213) );
  OAI2BB2X1 aes_core_keymem_U700 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[12]), .Y(aes_core_keymem_n2225) );
  OAI2BB2X1 aes_core_keymem_U699 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[11]), .Y(aes_core_keymem_n2237) );
  OAI2BB2X1 aes_core_keymem_U698 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[10]), .Y(aes_core_keymem_n2249) );
  OAI2BB2X1 aes_core_keymem_U697 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[9]), .Y(aes_core_keymem_n2261) );
  OAI2BB2X1 aes_core_keymem_U696 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[8]), .Y(aes_core_keymem_n2273) );
  OAI2BB2X1 aes_core_keymem_U695 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[7]), .Y(aes_core_keymem_n2285) );
  OAI2BB2X1 aes_core_keymem_U694 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[6]), .Y(aes_core_keymem_n2297) );
  OAI2BB2X1 aes_core_keymem_U693 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[5]), .Y(aes_core_keymem_n2309) );
  OAI2BB2X1 aes_core_keymem_U692 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[4]), .Y(aes_core_keymem_n2321) );
  OAI2BB2X1 aes_core_keymem_U691 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[3]), .Y(aes_core_keymem_n2333) );
  OAI2BB2X1 aes_core_keymem_U690 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[2]), .Y(aes_core_keymem_n2345) );
  OAI2BB2X1 aes_core_keymem_U689 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[1]), .Y(aes_core_keymem_n2357) );
  OAI2BB2X1 aes_core_keymem_U688 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n550), .A0N(aes_core_keymem_n550), .A1N(
        aes_core_keymem_key_mem[0]), .Y(aes_core_keymem_n2369) );
  OAI2BB2X1 aes_core_keymem_U687 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[383]), .Y(aes_core_keymem_n847) );
  OAI2BB2X1 aes_core_keymem_U686 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[382]), .Y(aes_core_keymem_n859) );
  OAI2BB2X1 aes_core_keymem_U685 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[381]), .Y(aes_core_keymem_n871) );
  OAI2BB2X1 aes_core_keymem_U684 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[380]), .Y(aes_core_keymem_n883) );
  OAI2BB2X1 aes_core_keymem_U683 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[379]), .Y(aes_core_keymem_n895) );
  OAI2BB2X1 aes_core_keymem_U682 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[378]), .Y(aes_core_keymem_n907) );
  OAI2BB2X1 aes_core_keymem_U681 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[377]), .Y(aes_core_keymem_n919) );
  OAI2BB2X1 aes_core_keymem_U680 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[376]), .Y(aes_core_keymem_n931) );
  OAI2BB2X1 aes_core_keymem_U679 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[375]), .Y(aes_core_keymem_n943) );
  OAI2BB2X1 aes_core_keymem_U678 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[374]), .Y(aes_core_keymem_n955) );
  OAI2BB2X1 aes_core_keymem_U677 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[373]), .Y(aes_core_keymem_n967) );
  OAI2BB2X1 aes_core_keymem_U676 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[372]), .Y(aes_core_keymem_n979) );
  OAI2BB2X1 aes_core_keymem_U675 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[371]), .Y(aes_core_keymem_n991) );
  OAI2BB2X1 aes_core_keymem_U674 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[370]), .Y(aes_core_keymem_n1003) );
  OAI2BB2X1 aes_core_keymem_U673 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[369]), .Y(aes_core_keymem_n1015) );
  OAI2BB2X1 aes_core_keymem_U672 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[368]), .Y(aes_core_keymem_n1027) );
  OAI2BB2X1 aes_core_keymem_U671 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[367]), .Y(aes_core_keymem_n1039) );
  OAI2BB2X1 aes_core_keymem_U670 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[366]), .Y(aes_core_keymem_n1051) );
  OAI2BB2X1 aes_core_keymem_U669 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[365]), .Y(aes_core_keymem_n1063) );
  OAI2BB2X1 aes_core_keymem_U668 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[364]), .Y(aes_core_keymem_n1075) );
  OAI2BB2X1 aes_core_keymem_U667 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[363]), .Y(aes_core_keymem_n1087) );
  OAI2BB2X1 aes_core_keymem_U666 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[362]), .Y(aes_core_keymem_n1099) );
  OAI2BB2X1 aes_core_keymem_U665 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[361]), .Y(aes_core_keymem_n1111) );
  OAI2BB2X1 aes_core_keymem_U664 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[360]), .Y(aes_core_keymem_n1123) );
  OAI2BB2X1 aes_core_keymem_U663 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[359]), .Y(aes_core_keymem_n1135) );
  OAI2BB2X1 aes_core_keymem_U662 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[358]), .Y(aes_core_keymem_n1147) );
  OAI2BB2X1 aes_core_keymem_U661 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[357]), .Y(aes_core_keymem_n1159) );
  OAI2BB2X1 aes_core_keymem_U660 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[356]), .Y(aes_core_keymem_n1171) );
  OAI2BB2X1 aes_core_keymem_U659 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[355]), .Y(aes_core_keymem_n1183) );
  OAI2BB2X1 aes_core_keymem_U658 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[354]), .Y(aes_core_keymem_n1195) );
  OAI2BB2X1 aes_core_keymem_U657 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[353]), .Y(aes_core_keymem_n1207) );
  OAI2BB2X1 aes_core_keymem_U656 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[352]), .Y(aes_core_keymem_n1219) );
  OAI2BB2X1 aes_core_keymem_U655 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[351]), .Y(aes_core_keymem_n1231) );
  OAI2BB2X1 aes_core_keymem_U654 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[350]), .Y(aes_core_keymem_n1243) );
  OAI2BB2X1 aes_core_keymem_U653 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[349]), .Y(aes_core_keymem_n1255) );
  OAI2BB2X1 aes_core_keymem_U652 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[348]), .Y(aes_core_keymem_n1267) );
  OAI2BB2X1 aes_core_keymem_U651 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[347]), .Y(aes_core_keymem_n1279) );
  OAI2BB2X1 aes_core_keymem_U650 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[346]), .Y(aes_core_keymem_n1291) );
  OAI2BB2X1 aes_core_keymem_U649 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[345]), .Y(aes_core_keymem_n1303) );
  OAI2BB2X1 aes_core_keymem_U648 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[344]), .Y(aes_core_keymem_n1315) );
  OAI2BB2X1 aes_core_keymem_U647 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[343]), .Y(aes_core_keymem_n1327) );
  OAI2BB2X1 aes_core_keymem_U646 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[342]), .Y(aes_core_keymem_n1339) );
  OAI2BB2X1 aes_core_keymem_U645 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[341]), .Y(aes_core_keymem_n1351) );
  OAI2BB2X1 aes_core_keymem_U644 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[340]), .Y(aes_core_keymem_n1363) );
  OAI2BB2X1 aes_core_keymem_U643 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[339]), .Y(aes_core_keymem_n1375) );
  OAI2BB2X1 aes_core_keymem_U642 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[338]), .Y(aes_core_keymem_n1387) );
  OAI2BB2X1 aes_core_keymem_U641 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[337]), .Y(aes_core_keymem_n1399) );
  OAI2BB2X1 aes_core_keymem_U640 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[336]), .Y(aes_core_keymem_n1411) );
  OAI2BB2X1 aes_core_keymem_U639 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[335]), .Y(aes_core_keymem_n1423) );
  OAI2BB2X1 aes_core_keymem_U638 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[334]), .Y(aes_core_keymem_n1435) );
  OAI2BB2X1 aes_core_keymem_U637 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[333]), .Y(aes_core_keymem_n1447) );
  OAI2BB2X1 aes_core_keymem_U636 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[332]), .Y(aes_core_keymem_n1459) );
  OAI2BB2X1 aes_core_keymem_U635 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[331]), .Y(aes_core_keymem_n1471) );
  OAI2BB2X1 aes_core_keymem_U634 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[330]), .Y(aes_core_keymem_n1483) );
  OAI2BB2X1 aes_core_keymem_U633 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[329]), .Y(aes_core_keymem_n1495) );
  OAI2BB2X1 aes_core_keymem_U632 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[328]), .Y(aes_core_keymem_n1507) );
  OAI2BB2X1 aes_core_keymem_U631 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[327]), .Y(aes_core_keymem_n1519) );
  OAI2BB2X1 aes_core_keymem_U630 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[326]), .Y(aes_core_keymem_n1531) );
  OAI2BB2X1 aes_core_keymem_U629 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[325]), .Y(aes_core_keymem_n1543) );
  OAI2BB2X1 aes_core_keymem_U628 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[324]), .Y(aes_core_keymem_n1555) );
  OAI2BB2X1 aes_core_keymem_U627 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[323]), .Y(aes_core_keymem_n1567) );
  OAI2BB2X1 aes_core_keymem_U626 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[322]), .Y(aes_core_keymem_n1579) );
  OAI2BB2X1 aes_core_keymem_U625 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[321]), .Y(aes_core_keymem_n1591) );
  OAI2BB2X1 aes_core_keymem_U624 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[320]), .Y(aes_core_keymem_n1603) );
  OAI2BB2X1 aes_core_keymem_U623 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[319]), .Y(aes_core_keymem_n1615) );
  OAI2BB2X1 aes_core_keymem_U622 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[318]), .Y(aes_core_keymem_n1627) );
  OAI2BB2X1 aes_core_keymem_U621 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[317]), .Y(aes_core_keymem_n1639) );
  OAI2BB2X1 aes_core_keymem_U620 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[316]), .Y(aes_core_keymem_n1651) );
  OAI2BB2X1 aes_core_keymem_U619 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[315]), .Y(aes_core_keymem_n1663) );
  OAI2BB2X1 aes_core_keymem_U618 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[314]), .Y(aes_core_keymem_n1675) );
  OAI2BB2X1 aes_core_keymem_U617 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[313]), .Y(aes_core_keymem_n1687) );
  OAI2BB2X1 aes_core_keymem_U616 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[312]), .Y(aes_core_keymem_n1699) );
  OAI2BB2X1 aes_core_keymem_U615 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[311]), .Y(aes_core_keymem_n1711) );
  OAI2BB2X1 aes_core_keymem_U614 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[310]), .Y(aes_core_keymem_n1723) );
  OAI2BB2X1 aes_core_keymem_U613 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[309]), .Y(aes_core_keymem_n1735) );
  OAI2BB2X1 aes_core_keymem_U612 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[308]), .Y(aes_core_keymem_n1747) );
  OAI2BB2X1 aes_core_keymem_U611 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[307]), .Y(aes_core_keymem_n1759) );
  OAI2BB2X1 aes_core_keymem_U610 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[306]), .Y(aes_core_keymem_n1771) );
  OAI2BB2X1 aes_core_keymem_U609 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[305]), .Y(aes_core_keymem_n1783) );
  OAI2BB2X1 aes_core_keymem_U608 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[304]), .Y(aes_core_keymem_n1795) );
  OAI2BB2X1 aes_core_keymem_U607 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[303]), .Y(aes_core_keymem_n1807) );
  OAI2BB2X1 aes_core_keymem_U606 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[302]), .Y(aes_core_keymem_n1819) );
  OAI2BB2X1 aes_core_keymem_U605 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[301]), .Y(aes_core_keymem_n1831) );
  OAI2BB2X1 aes_core_keymem_U604 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[300]), .Y(aes_core_keymem_n1843) );
  OAI2BB2X1 aes_core_keymem_U603 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[299]), .Y(aes_core_keymem_n1855) );
  OAI2BB2X1 aes_core_keymem_U602 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[298]), .Y(aes_core_keymem_n1867) );
  OAI2BB2X1 aes_core_keymem_U601 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[297]), .Y(aes_core_keymem_n1879) );
  OAI2BB2X1 aes_core_keymem_U600 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[296]), .Y(aes_core_keymem_n1891) );
  OAI2BB2X1 aes_core_keymem_U599 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[295]), .Y(aes_core_keymem_n1903) );
  OAI2BB2X1 aes_core_keymem_U598 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[294]), .Y(aes_core_keymem_n1915) );
  OAI2BB2X1 aes_core_keymem_U597 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[293]), .Y(aes_core_keymem_n1927) );
  OAI2BB2X1 aes_core_keymem_U596 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[292]), .Y(aes_core_keymem_n1939) );
  OAI2BB2X1 aes_core_keymem_U595 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[291]), .Y(aes_core_keymem_n1951) );
  OAI2BB2X1 aes_core_keymem_U594 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[290]), .Y(aes_core_keymem_n1963) );
  OAI2BB2X1 aes_core_keymem_U593 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[289]), .Y(aes_core_keymem_n1975) );
  OAI2BB2X1 aes_core_keymem_U592 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[288]), .Y(aes_core_keymem_n1987) );
  OAI2BB2X1 aes_core_keymem_U591 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[287]), .Y(aes_core_keymem_n1999) );
  OAI2BB2X1 aes_core_keymem_U590 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[286]), .Y(aes_core_keymem_n2011) );
  OAI2BB2X1 aes_core_keymem_U589 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[285]), .Y(aes_core_keymem_n2023) );
  OAI2BB2X1 aes_core_keymem_U588 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[284]), .Y(aes_core_keymem_n2035) );
  OAI2BB2X1 aes_core_keymem_U587 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[283]), .Y(aes_core_keymem_n2047) );
  OAI2BB2X1 aes_core_keymem_U586 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[282]), .Y(aes_core_keymem_n2059) );
  OAI2BB2X1 aes_core_keymem_U585 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[281]), .Y(aes_core_keymem_n2071) );
  OAI2BB2X1 aes_core_keymem_U584 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[280]), .Y(aes_core_keymem_n2083) );
  OAI2BB2X1 aes_core_keymem_U583 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[279]), .Y(aes_core_keymem_n2095) );
  OAI2BB2X1 aes_core_keymem_U582 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[278]), .Y(aes_core_keymem_n2107) );
  OAI2BB2X1 aes_core_keymem_U581 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[277]), .Y(aes_core_keymem_n2119) );
  OAI2BB2X1 aes_core_keymem_U580 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[276]), .Y(aes_core_keymem_n2131) );
  OAI2BB2X1 aes_core_keymem_U579 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[275]), .Y(aes_core_keymem_n2143) );
  OAI2BB2X1 aes_core_keymem_U578 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[274]), .Y(aes_core_keymem_n2155) );
  OAI2BB2X1 aes_core_keymem_U577 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[273]), .Y(aes_core_keymem_n2167) );
  OAI2BB2X1 aes_core_keymem_U576 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[272]), .Y(aes_core_keymem_n2179) );
  OAI2BB2X1 aes_core_keymem_U575 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[271]), .Y(aes_core_keymem_n2191) );
  OAI2BB2X1 aes_core_keymem_U574 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[270]), .Y(aes_core_keymem_n2203) );
  OAI2BB2X1 aes_core_keymem_U573 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[269]), .Y(aes_core_keymem_n2215) );
  OAI2BB2X1 aes_core_keymem_U572 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[268]), .Y(aes_core_keymem_n2227) );
  OAI2BB2X1 aes_core_keymem_U571 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[267]), .Y(aes_core_keymem_n2239) );
  OAI2BB2X1 aes_core_keymem_U570 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[266]), .Y(aes_core_keymem_n2251) );
  OAI2BB2X1 aes_core_keymem_U569 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[265]), .Y(aes_core_keymem_n2263) );
  OAI2BB2X1 aes_core_keymem_U568 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[264]), .Y(aes_core_keymem_n2275) );
  OAI2BB2X1 aes_core_keymem_U567 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[263]), .Y(aes_core_keymem_n2287) );
  OAI2BB2X1 aes_core_keymem_U566 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[262]), .Y(aes_core_keymem_n2299) );
  OAI2BB2X1 aes_core_keymem_U565 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[261]), .Y(aes_core_keymem_n2311) );
  OAI2BB2X1 aes_core_keymem_U564 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[260]), .Y(aes_core_keymem_n2323) );
  OAI2BB2X1 aes_core_keymem_U563 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[259]), .Y(aes_core_keymem_n2335) );
  OAI2BB2X1 aes_core_keymem_U562 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[258]), .Y(aes_core_keymem_n2347) );
  OAI2BB2X1 aes_core_keymem_U561 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[257]), .Y(aes_core_keymem_n2359) );
  OAI2BB2X1 aes_core_keymem_U560 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n552), .A0N(aes_core_keymem_n552), .A1N(
        aes_core_keymem_key_mem[256]), .Y(aes_core_keymem_n2371) );
  OAI2BB2X1 aes_core_keymem_U559 ( .B0(aes_core_keymem_n2505), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[639]), .Y(aes_core_keymem_n842) );
  OAI2BB2X1 aes_core_keymem_U558 ( .B0(aes_core_keymem_n2504), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[638]), .Y(aes_core_keymem_n854) );
  OAI2BB2X1 aes_core_keymem_U557 ( .B0(aes_core_keymem_n2503), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[637]), .Y(aes_core_keymem_n866) );
  OAI2BB2X1 aes_core_keymem_U556 ( .B0(aes_core_keymem_n2502), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[636]), .Y(aes_core_keymem_n878) );
  OAI2BB2X1 aes_core_keymem_U555 ( .B0(aes_core_keymem_n2501), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[635]), .Y(aes_core_keymem_n890) );
  OAI2BB2X1 aes_core_keymem_U554 ( .B0(aes_core_keymem_n2500), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[634]), .Y(aes_core_keymem_n902) );
  OAI2BB2X1 aes_core_keymem_U553 ( .B0(aes_core_keymem_n2499), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[633]), .Y(aes_core_keymem_n914) );
  OAI2BB2X1 aes_core_keymem_U552 ( .B0(aes_core_keymem_n2498), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[632]), .Y(aes_core_keymem_n926) );
  OAI2BB2X1 aes_core_keymem_U551 ( .B0(aes_core_keymem_n2497), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[631]), .Y(aes_core_keymem_n938) );
  OAI2BB2X1 aes_core_keymem_U550 ( .B0(aes_core_keymem_n2496), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[630]), .Y(aes_core_keymem_n950) );
  OAI2BB2X1 aes_core_keymem_U549 ( .B0(aes_core_keymem_n2495), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[629]), .Y(aes_core_keymem_n962) );
  OAI2BB2X1 aes_core_keymem_U548 ( .B0(aes_core_keymem_n2494), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[628]), .Y(aes_core_keymem_n974) );
  OAI2BB2X1 aes_core_keymem_U547 ( .B0(aes_core_keymem_n2493), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[627]), .Y(aes_core_keymem_n986) );
  OAI2BB2X1 aes_core_keymem_U546 ( .B0(aes_core_keymem_n2492), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[626]), .Y(aes_core_keymem_n998) );
  OAI2BB2X1 aes_core_keymem_U545 ( .B0(aes_core_keymem_n2491), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[625]), .Y(aes_core_keymem_n1010) );
  OAI2BB2X1 aes_core_keymem_U544 ( .B0(aes_core_keymem_n2490), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[624]), .Y(aes_core_keymem_n1022) );
  OAI2BB2X1 aes_core_keymem_U543 ( .B0(aes_core_keymem_n2489), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[623]), .Y(aes_core_keymem_n1034) );
  OAI2BB2X1 aes_core_keymem_U542 ( .B0(aes_core_keymem_n2488), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[622]), .Y(aes_core_keymem_n1046) );
  OAI2BB2X1 aes_core_keymem_U541 ( .B0(aes_core_keymem_n2487), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[621]), .Y(aes_core_keymem_n1058) );
  OAI2BB2X1 aes_core_keymem_U540 ( .B0(aes_core_keymem_n2486), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[620]), .Y(aes_core_keymem_n1070) );
  OAI2BB2X1 aes_core_keymem_U539 ( .B0(aes_core_keymem_n2485), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[619]), .Y(aes_core_keymem_n1082) );
  OAI2BB2X1 aes_core_keymem_U538 ( .B0(aes_core_keymem_n2484), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[618]), .Y(aes_core_keymem_n1094) );
  OAI2BB2X1 aes_core_keymem_U537 ( .B0(aes_core_keymem_n2483), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[617]), .Y(aes_core_keymem_n1106) );
  OAI2BB2X1 aes_core_keymem_U536 ( .B0(aes_core_keymem_n2482), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[616]), .Y(aes_core_keymem_n1118) );
  OAI2BB2X1 aes_core_keymem_U535 ( .B0(aes_core_keymem_n2481), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[615]), .Y(aes_core_keymem_n1130) );
  OAI2BB2X1 aes_core_keymem_U534 ( .B0(aes_core_keymem_n2480), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[614]), .Y(aes_core_keymem_n1142) );
  OAI2BB2X1 aes_core_keymem_U533 ( .B0(aes_core_keymem_n2479), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[613]), .Y(aes_core_keymem_n1154) );
  OAI2BB2X1 aes_core_keymem_U532 ( .B0(aes_core_keymem_n2478), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[612]), .Y(aes_core_keymem_n1166) );
  OAI2BB2X1 aes_core_keymem_U531 ( .B0(aes_core_keymem_n2477), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[611]), .Y(aes_core_keymem_n1178) );
  OAI2BB2X1 aes_core_keymem_U530 ( .B0(aes_core_keymem_n2476), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[610]), .Y(aes_core_keymem_n1190) );
  OAI2BB2X1 aes_core_keymem_U529 ( .B0(aes_core_keymem_n2475), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[609]), .Y(aes_core_keymem_n1202) );
  OAI2BB2X1 aes_core_keymem_U528 ( .B0(aes_core_keymem_n2474), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[608]), .Y(aes_core_keymem_n1214) );
  OAI2BB2X1 aes_core_keymem_U527 ( .B0(aes_core_keymem_n2473), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[607]), .Y(aes_core_keymem_n1226) );
  OAI2BB2X1 aes_core_keymem_U526 ( .B0(aes_core_keymem_n2472), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[606]), .Y(aes_core_keymem_n1238) );
  OAI2BB2X1 aes_core_keymem_U525 ( .B0(aes_core_keymem_n2471), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[605]), .Y(aes_core_keymem_n1250) );
  OAI2BB2X1 aes_core_keymem_U524 ( .B0(aes_core_keymem_n2470), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[604]), .Y(aes_core_keymem_n1262) );
  OAI2BB2X1 aes_core_keymem_U523 ( .B0(aes_core_keymem_n2469), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[603]), .Y(aes_core_keymem_n1274) );
  OAI2BB2X1 aes_core_keymem_U522 ( .B0(aes_core_keymem_n2468), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[602]), .Y(aes_core_keymem_n1286) );
  OAI2BB2X1 aes_core_keymem_U521 ( .B0(aes_core_keymem_n2467), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[601]), .Y(aes_core_keymem_n1298) );
  OAI2BB2X1 aes_core_keymem_U520 ( .B0(aes_core_keymem_n2466), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[600]), .Y(aes_core_keymem_n1310) );
  OAI2BB2X1 aes_core_keymem_U519 ( .B0(aes_core_keymem_n2465), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[599]), .Y(aes_core_keymem_n1322) );
  OAI2BB2X1 aes_core_keymem_U518 ( .B0(aes_core_keymem_n2464), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[598]), .Y(aes_core_keymem_n1334) );
  OAI2BB2X1 aes_core_keymem_U517 ( .B0(aes_core_keymem_n2463), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[597]), .Y(aes_core_keymem_n1346) );
  OAI2BB2X1 aes_core_keymem_U516 ( .B0(aes_core_keymem_n2462), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[596]), .Y(aes_core_keymem_n1358) );
  OAI2BB2X1 aes_core_keymem_U515 ( .B0(aes_core_keymem_n2461), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[595]), .Y(aes_core_keymem_n1370) );
  OAI2BB2X1 aes_core_keymem_U514 ( .B0(aes_core_keymem_n2460), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[594]), .Y(aes_core_keymem_n1382) );
  OAI2BB2X1 aes_core_keymem_U513 ( .B0(aes_core_keymem_n2459), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[593]), .Y(aes_core_keymem_n1394) );
  OAI2BB2X1 aes_core_keymem_U512 ( .B0(aes_core_keymem_n2458), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[592]), .Y(aes_core_keymem_n1406) );
  OAI2BB2X1 aes_core_keymem_U511 ( .B0(aes_core_keymem_n2457), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[591]), .Y(aes_core_keymem_n1418) );
  OAI2BB2X1 aes_core_keymem_U510 ( .B0(aes_core_keymem_n2456), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[590]), .Y(aes_core_keymem_n1430) );
  OAI2BB2X1 aes_core_keymem_U509 ( .B0(aes_core_keymem_n2455), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[589]), .Y(aes_core_keymem_n1442) );
  OAI2BB2X1 aes_core_keymem_U508 ( .B0(aes_core_keymem_n2454), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[588]), .Y(aes_core_keymem_n1454) );
  OAI2BB2X1 aes_core_keymem_U507 ( .B0(aes_core_keymem_n2453), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[587]), .Y(aes_core_keymem_n1466) );
  OAI2BB2X1 aes_core_keymem_U506 ( .B0(aes_core_keymem_n2452), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[586]), .Y(aes_core_keymem_n1478) );
  OAI2BB2X1 aes_core_keymem_U505 ( .B0(aes_core_keymem_n2451), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[585]), .Y(aes_core_keymem_n1490) );
  OAI2BB2X1 aes_core_keymem_U504 ( .B0(aes_core_keymem_n2450), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[584]), .Y(aes_core_keymem_n1502) );
  OAI2BB2X1 aes_core_keymem_U503 ( .B0(aes_core_keymem_n2449), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[583]), .Y(aes_core_keymem_n1514) );
  OAI2BB2X1 aes_core_keymem_U502 ( .B0(aes_core_keymem_n2448), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[582]), .Y(aes_core_keymem_n1526) );
  OAI2BB2X1 aes_core_keymem_U501 ( .B0(aes_core_keymem_n2447), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[581]), .Y(aes_core_keymem_n1538) );
  OAI2BB2X1 aes_core_keymem_U500 ( .B0(aes_core_keymem_n2446), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[580]), .Y(aes_core_keymem_n1550) );
  OAI2BB2X1 aes_core_keymem_U499 ( .B0(aes_core_keymem_n2445), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[579]), .Y(aes_core_keymem_n1562) );
  OAI2BB2X1 aes_core_keymem_U498 ( .B0(aes_core_keymem_n2444), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[578]), .Y(aes_core_keymem_n1574) );
  OAI2BB2X1 aes_core_keymem_U497 ( .B0(aes_core_keymem_n2443), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[577]), .Y(aes_core_keymem_n1586) );
  OAI2BB2X1 aes_core_keymem_U496 ( .B0(aes_core_keymem_n2442), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[576]), .Y(aes_core_keymem_n1598) );
  OAI2BB2X1 aes_core_keymem_U495 ( .B0(aes_core_keymem_n2441), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[575]), .Y(aes_core_keymem_n1610) );
  OAI2BB2X1 aes_core_keymem_U494 ( .B0(aes_core_keymem_n2440), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[574]), .Y(aes_core_keymem_n1622) );
  OAI2BB2X1 aes_core_keymem_U493 ( .B0(aes_core_keymem_n2439), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[573]), .Y(aes_core_keymem_n1634) );
  OAI2BB2X1 aes_core_keymem_U492 ( .B0(aes_core_keymem_n2438), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[572]), .Y(aes_core_keymem_n1646) );
  OAI2BB2X1 aes_core_keymem_U491 ( .B0(aes_core_keymem_n2437), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[571]), .Y(aes_core_keymem_n1658) );
  OAI2BB2X1 aes_core_keymem_U490 ( .B0(aes_core_keymem_n2436), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[570]), .Y(aes_core_keymem_n1670) );
  OAI2BB2X1 aes_core_keymem_U489 ( .B0(aes_core_keymem_n2435), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[569]), .Y(aes_core_keymem_n1682) );
  OAI2BB2X1 aes_core_keymem_U488 ( .B0(aes_core_keymem_n2434), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[568]), .Y(aes_core_keymem_n1694) );
  OAI2BB2X1 aes_core_keymem_U487 ( .B0(aes_core_keymem_n2433), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[567]), .Y(aes_core_keymem_n1706) );
  OAI2BB2X1 aes_core_keymem_U486 ( .B0(aes_core_keymem_n2432), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[566]), .Y(aes_core_keymem_n1718) );
  OAI2BB2X1 aes_core_keymem_U485 ( .B0(aes_core_keymem_n2431), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[565]), .Y(aes_core_keymem_n1730) );
  OAI2BB2X1 aes_core_keymem_U484 ( .B0(aes_core_keymem_n2430), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[564]), .Y(aes_core_keymem_n1742) );
  OAI2BB2X1 aes_core_keymem_U483 ( .B0(aes_core_keymem_n2429), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[563]), .Y(aes_core_keymem_n1754) );
  OAI2BB2X1 aes_core_keymem_U482 ( .B0(aes_core_keymem_n2428), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[562]), .Y(aes_core_keymem_n1766) );
  OAI2BB2X1 aes_core_keymem_U481 ( .B0(aes_core_keymem_n2427), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[561]), .Y(aes_core_keymem_n1778) );
  OAI2BB2X1 aes_core_keymem_U480 ( .B0(aes_core_keymem_n2426), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[560]), .Y(aes_core_keymem_n1790) );
  OAI2BB2X1 aes_core_keymem_U479 ( .B0(aes_core_keymem_n2425), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[559]), .Y(aes_core_keymem_n1802) );
  OAI2BB2X1 aes_core_keymem_U478 ( .B0(aes_core_keymem_n2424), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[558]), .Y(aes_core_keymem_n1814) );
  OAI2BB2X1 aes_core_keymem_U477 ( .B0(aes_core_keymem_n2423), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[557]), .Y(aes_core_keymem_n1826) );
  OAI2BB2X1 aes_core_keymem_U476 ( .B0(aes_core_keymem_n2422), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[556]), .Y(aes_core_keymem_n1838) );
  OAI2BB2X1 aes_core_keymem_U475 ( .B0(aes_core_keymem_n2421), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[555]), .Y(aes_core_keymem_n1850) );
  OAI2BB2X1 aes_core_keymem_U474 ( .B0(aes_core_keymem_n2420), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[554]), .Y(aes_core_keymem_n1862) );
  OAI2BB2X1 aes_core_keymem_U473 ( .B0(aes_core_keymem_n2419), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[553]), .Y(aes_core_keymem_n1874) );
  OAI2BB2X1 aes_core_keymem_U472 ( .B0(aes_core_keymem_n2418), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[552]), .Y(aes_core_keymem_n1886) );
  OAI2BB2X1 aes_core_keymem_U471 ( .B0(aes_core_keymem_n2417), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[551]), .Y(aes_core_keymem_n1898) );
  OAI2BB2X1 aes_core_keymem_U470 ( .B0(aes_core_keymem_n2416), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[550]), .Y(aes_core_keymem_n1910) );
  OAI2BB2X1 aes_core_keymem_U469 ( .B0(aes_core_keymem_n2415), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[549]), .Y(aes_core_keymem_n1922) );
  OAI2BB2X1 aes_core_keymem_U468 ( .B0(aes_core_keymem_n2414), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[548]), .Y(aes_core_keymem_n1934) );
  OAI2BB2X1 aes_core_keymem_U467 ( .B0(aes_core_keymem_n2413), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[547]), .Y(aes_core_keymem_n1946) );
  OAI2BB2X1 aes_core_keymem_U466 ( .B0(aes_core_keymem_n2412), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[546]), .Y(aes_core_keymem_n1958) );
  OAI2BB2X1 aes_core_keymem_U465 ( .B0(aes_core_keymem_n2411), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[545]), .Y(aes_core_keymem_n1970) );
  OAI2BB2X1 aes_core_keymem_U464 ( .B0(aes_core_keymem_n2410), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[544]), .Y(aes_core_keymem_n1982) );
  OAI2BB2X1 aes_core_keymem_U463 ( .B0(aes_core_keymem_n2409), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[543]), .Y(aes_core_keymem_n1994) );
  OAI2BB2X1 aes_core_keymem_U462 ( .B0(aes_core_keymem_n2408), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[542]), .Y(aes_core_keymem_n2006) );
  OAI2BB2X1 aes_core_keymem_U461 ( .B0(aes_core_keymem_n2407), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[541]), .Y(aes_core_keymem_n2018) );
  OAI2BB2X1 aes_core_keymem_U460 ( .B0(aes_core_keymem_n2406), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[540]), .Y(aes_core_keymem_n2030) );
  OAI2BB2X1 aes_core_keymem_U459 ( .B0(aes_core_keymem_n2405), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[539]), .Y(aes_core_keymem_n2042) );
  OAI2BB2X1 aes_core_keymem_U458 ( .B0(aes_core_keymem_n2404), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[538]), .Y(aes_core_keymem_n2054) );
  OAI2BB2X1 aes_core_keymem_U457 ( .B0(aes_core_keymem_n2403), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[537]), .Y(aes_core_keymem_n2066) );
  OAI2BB2X1 aes_core_keymem_U456 ( .B0(aes_core_keymem_n2402), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[536]), .Y(aes_core_keymem_n2078) );
  OAI2BB2X1 aes_core_keymem_U455 ( .B0(aes_core_keymem_n2401), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[535]), .Y(aes_core_keymem_n2090) );
  OAI2BB2X1 aes_core_keymem_U454 ( .B0(aes_core_keymem_n2400), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[534]), .Y(aes_core_keymem_n2102) );
  OAI2BB2X1 aes_core_keymem_U453 ( .B0(aes_core_keymem_n2399), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[533]), .Y(aes_core_keymem_n2114) );
  OAI2BB2X1 aes_core_keymem_U452 ( .B0(aes_core_keymem_n2398), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[532]), .Y(aes_core_keymem_n2126) );
  OAI2BB2X1 aes_core_keymem_U451 ( .B0(aes_core_keymem_n2397), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[531]), .Y(aes_core_keymem_n2138) );
  OAI2BB2X1 aes_core_keymem_U450 ( .B0(aes_core_keymem_n2396), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[530]), .Y(aes_core_keymem_n2150) );
  OAI2BB2X1 aes_core_keymem_U449 ( .B0(aes_core_keymem_n2395), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[529]), .Y(aes_core_keymem_n2162) );
  OAI2BB2X1 aes_core_keymem_U448 ( .B0(aes_core_keymem_n2394), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[528]), .Y(aes_core_keymem_n2174) );
  OAI2BB2X1 aes_core_keymem_U447 ( .B0(aes_core_keymem_n2393), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[527]), .Y(aes_core_keymem_n2186) );
  OAI2BB2X1 aes_core_keymem_U446 ( .B0(aes_core_keymem_n2392), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[526]), .Y(aes_core_keymem_n2198) );
  OAI2BB2X1 aes_core_keymem_U445 ( .B0(aes_core_keymem_n2391), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[525]), .Y(aes_core_keymem_n2210) );
  OAI2BB2X1 aes_core_keymem_U444 ( .B0(aes_core_keymem_n773), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[524]), .Y(aes_core_keymem_n2222) );
  OAI2BB2X1 aes_core_keymem_U443 ( .B0(aes_core_keymem_n770), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[523]), .Y(aes_core_keymem_n2234) );
  OAI2BB2X1 aes_core_keymem_U442 ( .B0(aes_core_keymem_n767), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[522]), .Y(aes_core_keymem_n2246) );
  OAI2BB2X1 aes_core_keymem_U441 ( .B0(aes_core_keymem_n764), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[521]), .Y(aes_core_keymem_n2258) );
  OAI2BB2X1 aes_core_keymem_U440 ( .B0(aes_core_keymem_n761), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[520]), .Y(aes_core_keymem_n2270) );
  OAI2BB2X1 aes_core_keymem_U439 ( .B0(aes_core_keymem_n758), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[519]), .Y(aes_core_keymem_n2282) );
  OAI2BB2X1 aes_core_keymem_U438 ( .B0(aes_core_keymem_n755), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[518]), .Y(aes_core_keymem_n2294) );
  OAI2BB2X1 aes_core_keymem_U437 ( .B0(aes_core_keymem_n752), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[517]), .Y(aes_core_keymem_n2306) );
  OAI2BB2X1 aes_core_keymem_U436 ( .B0(aes_core_keymem_n559), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[516]), .Y(aes_core_keymem_n2318) );
  OAI2BB2X1 aes_core_keymem_U435 ( .B0(aes_core_keymem_n557), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[515]), .Y(aes_core_keymem_n2330) );
  OAI2BB2X1 aes_core_keymem_U434 ( .B0(aes_core_keymem_n554), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[514]), .Y(aes_core_keymem_n2342) );
  OAI2BB2X1 aes_core_keymem_U433 ( .B0(aes_core_keymem_n544), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[513]), .Y(aes_core_keymem_n2354) );
  OAI2BB2X1 aes_core_keymem_U432 ( .B0(aes_core_keymem_n30), .B1(
        aes_core_keymem_n547), .A0N(aes_core_keymem_n547), .A1N(
        aes_core_keymem_key_mem[512]), .Y(aes_core_keymem_n2366) );
  OAI211X1 aes_core_keymem_U431 ( .A0(aes_core_keymem_n840), .A1(
        aes_core_keymem_n2765), .B0(aes_core_keymem_n838), .C0(
        aes_core_keymem_n829), .Y(aes_core_keymem_n2388) );
  OAI221X1 aes_core_keymem_U430 ( .A0(aes_core_keymem_n829), .A1(
        aes_core_keymem_n821), .B0(aes_core_keymem_n840), .B1(
        aes_core_keymem_n17), .C0(aes_core_keymem_n545), .Y(
        aes_core_keymem_n2390) );
  INVX1 aes_core_keymem_U429 ( .A(aes_core_keymem_n26), .Y(
        aes_core_keymem_n2716) );
  INVX1 aes_core_keymem_U428 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2728) );
  INVX1 aes_core_keymem_U427 ( .A(aes_core_keymem_n23), .Y(
        aes_core_keymem_n2749) );
  INVX1 aes_core_keymem_U426 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2739) );
  INVX1 aes_core_keymem_U425 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2706) );
  AOI21X1 aes_core_keymem_U424 ( .A0(aes_core_keymem_n2762), .A1(
        aes_core_keymem_n2768), .B0(aes_core_keymem_n836), .Y(
        aes_core_keymem_n837) );
  INVX1 aes_core_keymem_U423 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2750) );
  INVX1 aes_core_keymem_U422 ( .A(aes_core_keymem_n27), .Y(
        aes_core_keymem_n2705) );
  INVX1 aes_core_keymem_U421 ( .A(aes_core_keymem_n25), .Y(
        aes_core_keymem_n2727) );
  INVX1 aes_core_keymem_U420 ( .A(aes_core_keymem_n29), .Y(
        aes_core_keymem_n2683) );
  INVX1 aes_core_keymem_U419 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2662) );
  INVX1 aes_core_keymem_U418 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2695) );
  INVX1 aes_core_keymem_U417 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2673) );
  INVX1 aes_core_keymem_U416 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2717) );
  INVX1 aes_core_keymem_U415 ( .A(aes_core_keymem_n28), .Y(
        aes_core_keymem_n2694) );
  INVX1 aes_core_keymem_U414 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2684) );
  AOI32X1 aes_core_keymem_U413 ( .A0(aes_core_keymem_n825), .A1(
        aes_core_keymem_n2762), .A2(aes_core_keymem_n826), .B0(
        aes_core_keymem_n823), .B1(aes_core_keymem_n2762), .Y(
        aes_core_keymem_n839) );
  OAI21X1 aes_core_keymem_U412 ( .A0(aes_core_keymem_n837), .A1(
        aes_core_keymem_n2764), .B0(aes_core_keymem_n839), .Y(
        aes_core_keymem_n2389) );
  INVX1 aes_core_keymem_U411 ( .A(aes_core_keymem_n31), .Y(
        aes_core_keymem_n2661) );
  INVX1 aes_core_keymem_U410 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2652) );
  NAND3X1 aes_core_keymem_U409 ( .A(aes_core_keymem_n2762), .B(
        aes_core_keymem_n828), .C(aes_core_keymem_n827), .Y(
        aes_core_keymem_n555) );
  NAND3X1 aes_core_keymem_U408 ( .A(aes_core_keymem_n2762), .B(
        aes_core_keymem_n828), .C(aes_core_keymem_n824), .Y(
        aes_core_keymem_n556) );
  AND2X2 aes_core_keymem_U407 ( .A(aes_core_keymem_n542), .B(
        aes_core_keymem_n541), .Y(aes_core_keymem_n32) );
  NAND2X1 aes_core_keymem_U406 ( .A(aes_core_keymem_n823), .B(
        aes_core_keymem_n827), .Y(aes_core_keymem_n821) );
  NOR2X1 aes_core_keymem_U405 ( .A(aes_core_keymem_n2767), .B(
        aes_core_keymem_n2768), .Y(aes_core_keymem_n825) );
  INVX1 aes_core_keymem_U404 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2581) );
  INVX1 aes_core_keymem_U403 ( .A(aes_core_keymem_n17), .Y(aes_core_keymem_n24) );
  INVX1 aes_core_keymem_U402 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2738) );
  INVX1 aes_core_keymem_U401 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2715) );
  INVX1 aes_core_keymem_U400 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2730) );
  INVX1 aes_core_keymem_U399 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2732) );
  INVX1 aes_core_keymem_U398 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2735) );
  INVX1 aes_core_keymem_U397 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2737) );
  INVX1 aes_core_keymem_U396 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2731) );
  INVX1 aes_core_keymem_U395 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2734) );
  INVX1 aes_core_keymem_U394 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2733) );
  INVX1 aes_core_keymem_U393 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2729) );
  INVX1 aes_core_keymem_U392 ( .A(aes_core_keymem_n5), .Y(
        aes_core_keymem_n2736) );
  INVX1 aes_core_keymem_U391 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2741) );
  INVX1 aes_core_keymem_U390 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2743) );
  INVX1 aes_core_keymem_U389 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2709) );
  INVX1 aes_core_keymem_U388 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2746) );
  INVX1 aes_core_keymem_U387 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2712) );
  INVX1 aes_core_keymem_U386 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2748) );
  INVX1 aes_core_keymem_U385 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2714) );
  INVX1 aes_core_keymem_U384 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2742) );
  INVX1 aes_core_keymem_U383 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2708) );
  INVX1 aes_core_keymem_U382 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2745) );
  INVX1 aes_core_keymem_U381 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2711) );
  INVX1 aes_core_keymem_U380 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2744) );
  INVX1 aes_core_keymem_U379 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2710) );
  INVX1 aes_core_keymem_U378 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2740) );
  INVX1 aes_core_keymem_U377 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2707) );
  INVX1 aes_core_keymem_U376 ( .A(aes_core_keymem_n2749), .Y(
        aes_core_keymem_n2747) );
  INVX1 aes_core_keymem_U375 ( .A(aes_core_keymem_n2716), .Y(
        aes_core_keymem_n2713) );
  NAND2X1 aes_core_keymem_U374 ( .A(aes_core_keymem_n838), .B(
        aes_core_keymem_n829), .Y(aes_core_keymem_n834) );
  INVX1 aes_core_keymem_U373 ( .A(aes_core_keymem_n32), .Y(
        aes_core_keymem_n2651) );
  INVX1 aes_core_keymem_U372 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2704) );
  INVX1 aes_core_keymem_U371 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2682) );
  INVX1 aes_core_keymem_U370 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2760) );
  INVX1 aes_core_keymem_U369 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2726) );
  INVX1 aes_core_keymem_U368 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2697) );
  INVX1 aes_core_keymem_U367 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2699) );
  INVX1 aes_core_keymem_U366 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2703) );
  INVX1 aes_core_keymem_U365 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2698) );
  INVX1 aes_core_keymem_U364 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2701) );
  INVX1 aes_core_keymem_U363 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2700) );
  INVX1 aes_core_keymem_U362 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2663) );
  INVX1 aes_core_keymem_U361 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2696) );
  INVX1 aes_core_keymem_U360 ( .A(aes_core_keymem_n2705), .Y(
        aes_core_keymem_n2702) );
  INVX1 aes_core_keymem_U359 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2681) );
  INVX1 aes_core_keymem_U358 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2675) );
  INVX1 aes_core_keymem_U357 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2679) );
  INVX1 aes_core_keymem_U356 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2677) );
  INVX1 aes_core_keymem_U355 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2676) );
  INVX1 aes_core_keymem_U354 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2678) );
  INVX1 aes_core_keymem_U353 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2680) );
  INVX1 aes_core_keymem_U352 ( .A(aes_core_keymem_n2683), .Y(
        aes_core_keymem_n2674) );
  INVX1 aes_core_keymem_U351 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2752) );
  INVX1 aes_core_keymem_U350 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2719) );
  INVX1 aes_core_keymem_U349 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2754) );
  INVX1 aes_core_keymem_U348 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2757) );
  INVX1 aes_core_keymem_U347 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2723) );
  INVX1 aes_core_keymem_U346 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2759) );
  INVX1 aes_core_keymem_U345 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2725) );
  INVX1 aes_core_keymem_U344 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2693) );
  INVX1 aes_core_keymem_U343 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2753) );
  INVX1 aes_core_keymem_U342 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2720) );
  INVX1 aes_core_keymem_U341 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2687) );
  INVX1 aes_core_keymem_U340 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2756) );
  INVX1 aes_core_keymem_U339 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2722) );
  INVX1 aes_core_keymem_U338 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2691) );
  INVX1 aes_core_keymem_U337 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2755) );
  INVX1 aes_core_keymem_U336 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2721) );
  INVX1 aes_core_keymem_U335 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2689) );
  INVX1 aes_core_keymem_U334 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2688) );
  INVX1 aes_core_keymem_U333 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2690) );
  INVX1 aes_core_keymem_U332 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2751) );
  INVX1 aes_core_keymem_U331 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2718) );
  INVX1 aes_core_keymem_U330 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2686) );
  INVX1 aes_core_keymem_U329 ( .A(aes_core_keymem_n4), .Y(
        aes_core_keymem_n2758) );
  INVX1 aes_core_keymem_U328 ( .A(aes_core_keymem_n2727), .Y(
        aes_core_keymem_n2724) );
  INVX1 aes_core_keymem_U327 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2692) );
  INVX1 aes_core_keymem_U326 ( .A(aes_core_keymem_n2694), .Y(
        aes_core_keymem_n2685) );
  INVX1 aes_core_keymem_U325 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2642) );
  INVX1 aes_core_keymem_U324 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2655) );
  INVX1 aes_core_keymem_U323 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2658) );
  INVX1 aes_core_keymem_U322 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2660) );
  INVX1 aes_core_keymem_U321 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2654) );
  INVX1 aes_core_keymem_U320 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2657) );
  INVX1 aes_core_keymem_U319 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2656) );
  INVX1 aes_core_keymem_U318 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2653) );
  INVX1 aes_core_keymem_U317 ( .A(aes_core_keymem_n2661), .Y(
        aes_core_keymem_n2659) );
  INVX1 aes_core_keymem_U316 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2582) );
  INVX1 aes_core_keymem_U315 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2583) );
  INVX1 aes_core_keymem_U314 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2584) );
  INVX1 aes_core_keymem_U313 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2585) );
  INVX1 aes_core_keymem_U312 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2586) );
  INVX1 aes_core_keymem_U311 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2587) );
  INVX1 aes_core_keymem_U310 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2588) );
  INVX1 aes_core_keymem_U309 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2589) );
  INVX1 aes_core_keymem_U308 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2590) );
  INVX1 aes_core_keymem_U307 ( .A(aes_core_keymem_n1), .Y(
        aes_core_keymem_n2580) );
  INVX1 aes_core_keymem_U306 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2609) );
  INVX1 aes_core_keymem_U305 ( .A(aes_core_keymem_n3), .Y(
        aes_core_keymem_n2591) );
  INVX1 aes_core_keymem_U304 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2672) );
  INVX1 aes_core_keymem_U303 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2666) );
  INVX1 aes_core_keymem_U302 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2670) );
  INVX1 aes_core_keymem_U301 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2668) );
  INVX1 aes_core_keymem_U300 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2667) );
  INVX1 aes_core_keymem_U299 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2669) );
  INVX1 aes_core_keymem_U298 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2665) );
  INVX1 aes_core_keymem_U297 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2671) );
  INVX1 aes_core_keymem_U296 ( .A(aes_core_keymem_n16), .Y(
        aes_core_keymem_n2664) );
  INVX1 aes_core_keymem_U295 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2644) );
  INVX1 aes_core_keymem_U294 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2648) );
  INVX1 aes_core_keymem_U293 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2650) );
  INVX1 aes_core_keymem_U292 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2645) );
  INVX1 aes_core_keymem_U291 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2647) );
  INVX1 aes_core_keymem_U290 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2646) );
  INVX1 aes_core_keymem_U289 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2643) );
  INVX1 aes_core_keymem_U288 ( .A(aes_core_keymem_n2651), .Y(
        aes_core_keymem_n2649) );
  INVX1 aes_core_keymem_U287 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2626) );
  INVX1 aes_core_keymem_U286 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2610) );
  INVX1 aes_core_keymem_U285 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2592) );
  INVX1 aes_core_keymem_U284 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2593) );
  INVX1 aes_core_keymem_U283 ( .A(aes_core_keymem_n2638), .Y(
        aes_core_keymem_n2641) );
  INVX1 aes_core_keymem_U282 ( .A(aes_core_keymem_n2580), .Y(
        aes_core_keymem_n2574) );
  INVX1 aes_core_keymem_U281 ( .A(aes_core_keymem_n2556), .Y(
        aes_core_keymem_n2575) );
  INVX1 aes_core_keymem_U280 ( .A(aes_core_keymem_n2580), .Y(
        aes_core_keymem_n2576) );
  INVX1 aes_core_keymem_U279 ( .A(aes_core_keymem_n2580), .Y(
        aes_core_keymem_n2577) );
  INVX1 aes_core_keymem_U278 ( .A(aes_core_keymem_n2556), .Y(
        aes_core_keymem_n2578) );
  INVX1 aes_core_keymem_U277 ( .A(aes_core_keymem_n2556), .Y(
        aes_core_keymem_n2579) );
  INVX1 aes_core_keymem_U276 ( .A(aes_core_keymem_n2574), .Y(
        aes_core_keymem_n2573) );
  INVX1 aes_core_keymem_U275 ( .A(aes_core_keymem_n2573), .Y(
        aes_core_keymem_n2522) );
  INVX1 aes_core_keymem_U274 ( .A(aes_core_keymem_n2574), .Y(
        aes_core_keymem_n2572) );
  INVX1 aes_core_keymem_U273 ( .A(aes_core_keymem_n2574), .Y(
        aes_core_keymem_n2571) );
  INVX1 aes_core_keymem_U272 ( .A(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n2570) );
  INVX1 aes_core_keymem_U271 ( .A(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n2569) );
  INVX1 aes_core_keymem_U270 ( .A(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n2568) );
  INVX1 aes_core_keymem_U269 ( .A(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n2567) );
  INVX1 aes_core_keymem_U268 ( .A(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n2566) );
  INVX1 aes_core_keymem_U267 ( .A(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n2565) );
  INVX1 aes_core_keymem_U266 ( .A(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n2564) );
  INVX1 aes_core_keymem_U265 ( .A(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n2563) );
  INVX1 aes_core_keymem_U264 ( .A(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n2562) );
  INVX1 aes_core_keymem_U263 ( .A(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n2561) );
  INVX1 aes_core_keymem_U262 ( .A(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n2560) );
  INVX1 aes_core_keymem_U261 ( .A(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n2559) );
  INVX1 aes_core_keymem_U260 ( .A(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n2558) );
  INVX1 aes_core_keymem_U259 ( .A(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n2557) );
  INVX1 aes_core_keymem_U258 ( .A(aes_core_keymem_n1), .Y(
        aes_core_keymem_n2556) );
  INVX1 aes_core_keymem_U257 ( .A(aes_core_keymem_n2574), .Y(
        aes_core_keymem_n2555) );
  INVX1 aes_core_keymem_U256 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2615) );
  INVX1 aes_core_keymem_U255 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2598) );
  INVX1 aes_core_keymem_U254 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2627) );
  INVX1 aes_core_keymem_U253 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2611) );
  INVX1 aes_core_keymem_U252 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2594) );
  INVX1 aes_core_keymem_U251 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2628) );
  INVX1 aes_core_keymem_U250 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2612) );
  INVX1 aes_core_keymem_U249 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2595) );
  INVX1 aes_core_keymem_U248 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2629) );
  INVX1 aes_core_keymem_U247 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2613) );
  INVX1 aes_core_keymem_U246 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2596) );
  INVX1 aes_core_keymem_U245 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2630) );
  INVX1 aes_core_keymem_U244 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2614) );
  INVX1 aes_core_keymem_U243 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2597) );
  INVX1 aes_core_keymem_U242 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2617) );
  INVX1 aes_core_keymem_U241 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2600) );
  INVX1 aes_core_keymem_U240 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2616) );
  INVX1 aes_core_keymem_U239 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2599) );
  INVX1 aes_core_keymem_U238 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2633) );
  INVX1 aes_core_keymem_U237 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2618) );
  INVX1 aes_core_keymem_U236 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2601) );
  INVX1 aes_core_keymem_U235 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2619) );
  INVX1 aes_core_keymem_U234 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2602) );
  CLKINVX3 aes_core_keymem_U233 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2635) );
  CLKINVX3 aes_core_keymem_U232 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2620) );
  CLKINVX3 aes_core_keymem_U231 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2603) );
  CLKINVX3 aes_core_keymem_U230 ( .A(aes_core_keymem_n2641), .Y(
        aes_core_keymem_n2636) );
  CLKINVX3 aes_core_keymem_U229 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2637) );
  CLKINVX3 aes_core_keymem_U228 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2638) );
  CLKINVX3 aes_core_keymem_U227 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2621) );
  CLKINVX3 aes_core_keymem_U226 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2604) );
  CLKINVX3 aes_core_keymem_U225 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2639) );
  CLKINVX3 aes_core_keymem_U224 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2622) );
  CLKINVX3 aes_core_keymem_U223 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2605) );
  CLKINVX3 aes_core_keymem_U222 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2640) );
  CLKINVX3 aes_core_keymem_U221 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2623) );
  CLKINVX3 aes_core_keymem_U220 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2606) );
  CLKINVX3 aes_core_keymem_U219 ( .A(aes_core_keymem_n2625), .Y(
        aes_core_keymem_n2624) );
  CLKINVX3 aes_core_keymem_U218 ( .A(aes_core_keymem_n2608), .Y(
        aes_core_keymem_n2607) );
  INVX1 aes_core_keymem_U217 ( .A(aes_core_keymem_n2556), .Y(
        aes_core_keymem_n2554) );
  INVX1 aes_core_keymem_U216 ( .A(aes_core_keymem_n2572), .Y(
        aes_core_keymem_n2523) );
  INVX1 aes_core_keymem_U215 ( .A(aes_core_keymem_n2572), .Y(
        aes_core_keymem_n2524) );
  INVX1 aes_core_keymem_U214 ( .A(aes_core_keymem_n2571), .Y(
        aes_core_keymem_n2525) );
  INVX1 aes_core_keymem_U213 ( .A(aes_core_keymem_n2571), .Y(
        aes_core_keymem_n2526) );
  INVX1 aes_core_keymem_U212 ( .A(aes_core_keymem_n2570), .Y(
        aes_core_keymem_n2527) );
  INVX1 aes_core_keymem_U211 ( .A(aes_core_keymem_n2570), .Y(
        aes_core_keymem_n2528) );
  INVX1 aes_core_keymem_U210 ( .A(aes_core_keymem_n2569), .Y(
        aes_core_keymem_n2529) );
  INVX1 aes_core_keymem_U209 ( .A(aes_core_keymem_n2569), .Y(
        aes_core_keymem_n2530) );
  INVX1 aes_core_keymem_U208 ( .A(aes_core_keymem_n2568), .Y(
        aes_core_keymem_n2531) );
  INVX1 aes_core_keymem_U207 ( .A(aes_core_keymem_n2567), .Y(
        aes_core_keymem_n2532) );
  INVX1 aes_core_keymem_U206 ( .A(aes_core_keymem_n2567), .Y(
        aes_core_keymem_n2533) );
  INVX1 aes_core_keymem_U205 ( .A(aes_core_keymem_n2566), .Y(
        aes_core_keymem_n2534) );
  INVX1 aes_core_keymem_U204 ( .A(aes_core_keymem_n2566), .Y(
        aes_core_keymem_n2535) );
  INVX1 aes_core_keymem_U203 ( .A(aes_core_keymem_n2565), .Y(
        aes_core_keymem_n2536) );
  INVX1 aes_core_keymem_U202 ( .A(aes_core_keymem_n2565), .Y(
        aes_core_keymem_n2537) );
  INVX1 aes_core_keymem_U201 ( .A(aes_core_keymem_n2564), .Y(
        aes_core_keymem_n2538) );
  INVX1 aes_core_keymem_U200 ( .A(aes_core_keymem_n2563), .Y(
        aes_core_keymem_n2539) );
  INVX1 aes_core_keymem_U199 ( .A(aes_core_keymem_n2563), .Y(
        aes_core_keymem_n2540) );
  INVX1 aes_core_keymem_U198 ( .A(aes_core_keymem_n2562), .Y(
        aes_core_keymem_n2541) );
  INVX1 aes_core_keymem_U197 ( .A(aes_core_keymem_n2561), .Y(
        aes_core_keymem_n2542) );
  INVX1 aes_core_keymem_U196 ( .A(aes_core_keymem_n2561), .Y(
        aes_core_keymem_n2543) );
  INVX1 aes_core_keymem_U195 ( .A(aes_core_keymem_n2560), .Y(
        aes_core_keymem_n2544) );
  INVX1 aes_core_keymem_U194 ( .A(aes_core_keymem_n2560), .Y(
        aes_core_keymem_n2545) );
  INVX1 aes_core_keymem_U193 ( .A(aes_core_keymem_n2559), .Y(
        aes_core_keymem_n2546) );
  INVX1 aes_core_keymem_U192 ( .A(aes_core_keymem_n2559), .Y(
        aes_core_keymem_n2547) );
  INVX1 aes_core_keymem_U191 ( .A(aes_core_keymem_n2558), .Y(
        aes_core_keymem_n2548) );
  INVX1 aes_core_keymem_U190 ( .A(aes_core_keymem_n2557), .Y(
        aes_core_keymem_n2549) );
  INVX1 aes_core_keymem_U189 ( .A(aes_core_keymem_n2555), .Y(
        aes_core_keymem_n2551) );
  INVX1 aes_core_keymem_U188 ( .A(aes_core_keymem_n2573), .Y(
        aes_core_keymem_n2552) );
  INVX1 aes_core_keymem_U187 ( .A(aes_core_keymem_n2580), .Y(
        aes_core_keymem_n2553) );
  INVX1 aes_core_keymem_U186 ( .A(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n2511) );
  INVX1 aes_core_keymem_U185 ( .A(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n2506) );
  INVX1 aes_core_keymem_U184 ( .A(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n2507) );
  INVX1 aes_core_keymem_U183 ( .A(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n2508) );
  INVX1 aes_core_keymem_U182 ( .A(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n2509) );
  INVX1 aes_core_keymem_U181 ( .A(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n2510) );
  INVX1 aes_core_keymem_U180 ( .A(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n2513) );
  INVX1 aes_core_keymem_U179 ( .A(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n2512) );
  INVX1 aes_core_keymem_U178 ( .A(aes_core_keymem_n2576), .Y(
        aes_core_keymem_n2514) );
  INVX1 aes_core_keymem_U177 ( .A(aes_core_keymem_n2579), .Y(
        aes_core_keymem_n2515) );
  CLKINVX3 aes_core_keymem_U176 ( .A(aes_core_keymem_n2575), .Y(
        aes_core_keymem_n2516) );
  CLKINVX3 aes_core_keymem_U175 ( .A(aes_core_keymem_n2554), .Y(
        aes_core_keymem_n2517) );
  CLKINVX3 aes_core_keymem_U174 ( .A(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n2518) );
  CLKINVX3 aes_core_keymem_U173 ( .A(aes_core_keymem_n2577), .Y(
        aes_core_keymem_n2519) );
  CLKINVX3 aes_core_keymem_U172 ( .A(aes_core_keymem_n1), .Y(
        aes_core_keymem_n2520) );
  CLKINVX3 aes_core_keymem_U171 ( .A(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n2521) );
  AND3X1 aes_core_keymem_U170 ( .A(aes_core_enc_round_nr[1]), .B(
        aes_core_keymem_n2771), .C(aes_core_keymem_n542), .Y(
        aes_core_keymem_n28) );
  AND3X1 aes_core_keymem_U169 ( .A(aes_core_enc_round_nr[1]), .B(
        aes_core_keymem_n2771), .C(aes_core_enc_round_nr[2]), .Y(
        aes_core_keymem_n27) );
  AND3X1 aes_core_keymem_U168 ( .A(aes_core_enc_round_nr[0]), .B(
        aes_core_keymem_n2772), .C(aes_core_enc_round_nr[2]), .Y(
        aes_core_keymem_n25) );
  AND2X1 aes_core_keymem_U167 ( .A(aes_core_enc_round_nr[2]), .B(
        aes_core_keymem_n541), .Y(aes_core_keymem_n29) );
  OR3X1 aes_core_keymem_U166 ( .A(aes_core_keymem_n2772), .B(
        aes_core_enc_round_nr[2]), .C(aes_core_keymem_n2771), .Y(
        aes_core_keymem_n16) );
  INVX1 aes_core_keymem_U165 ( .A(aes_core_keymem_round_ctr_reg[3]), .Y(
        aes_core_keymem_n2764) );
  INVX1 aes_core_keymem_U164 ( .A(aes_core_keymem_round_ctr_reg[2]), .Y(
        aes_core_keymem_n2769) );
  NOR2X1 aes_core_keymem_U163 ( .A(aes_core_keymem_n2768), .B(
        aes_core_keymem_round_ctr_reg[0]), .Y(aes_core_keymem_n827) );
  AOI22X4 aes_core_keymem_U162 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n819), .B0(Din[129]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n818) );
  XOR2X2 aes_core_keymem_U161 ( .A(aes_core_keymem_prev_key1_reg[98]), .B(
        aes_core_new_sboxw[26]), .Y(aes_core_keymem_n617) );
  XOR2X2 aes_core_keymem_U160 ( .A(aes_core_keymem_prev_key1_reg[101]), .B(
        aes_core_new_sboxw[29]), .Y(aes_core_keymem_n611) );
  XOR2X2 aes_core_keymem_U159 ( .A(aes_core_keymem_prev_key1_reg[102]), .B(
        aes_core_new_sboxw[30]), .Y(aes_core_keymem_n609) );
  XOR2X1 aes_core_keymem_U158 ( .A(aes_core_keymem_prev_key1_reg[122]), .B(
        aes_core_keymem_rcon_reg[2]), .Y(aes_core_keymem_n15) );
  XOR2X1 aes_core_keymem_U157 ( .A(aes_core_keymem_prev_key1_reg[123]), .B(
        aes_core_keymem_rcon_reg[3]), .Y(aes_core_keymem_n13) );
  XOR2X1 aes_core_keymem_U156 ( .A(aes_core_keymem_prev_key1_reg[120]), .B(
        aes_core_keymem_rcon_reg[0]), .Y(aes_core_keymem_n12) );
  XOR2X1 aes_core_keymem_U155 ( .A(aes_core_keymem_prev_key1_reg[121]), .B(
        aes_core_keymem_rcon_reg[1]), .Y(aes_core_keymem_n11) );
  XOR2X1 aes_core_keymem_U154 ( .A(aes_core_keymem_prev_key1_reg[125]), .B(
        aes_core_keymem_rcon_reg[5]), .Y(aes_core_keymem_n10) );
  AOI22X4 aes_core_keymem_U153 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n809), .B0(Din[134]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n808) );
  AOI22X2 aes_core_keymem_U152 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n807), .B0(Din[135]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n806) );
  XOR2X2 aes_core_keymem_U151 ( .A(aes_core_keymem_n721), .B(
        aes_core_keymem_sboxw[14]), .Y(aes_core_keymem_n793) );
  BUFX12 aes_core_keymem_U150 ( .A(aes_core_keymem_n792), .Y(
        aes_core_keymem_n2392) );
  AOI22X2 aes_core_keymem_U149 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n769), .B0(Din[153]), .B1(aes_core_keymem_n2524), .Y(
        aes_core_keymem_n768) );
  XOR2X2 aes_core_keymem_U148 ( .A(aes_core_keymem_n723), .B(
        aes_core_keymem_sboxw[13]), .Y(aes_core_keymem_n795) );
  BUFX12 aes_core_keymem_U147 ( .A(aes_core_keymem_n794), .Y(
        aes_core_keymem_n2391) );
  AOI22X2 aes_core_keymem_U146 ( .A0(aes_core_keymem_n2589), .A1(
        aes_core_keymem_n766), .B0(Din[154]), .B1(aes_core_keymem_n2523), .Y(
        aes_core_keymem_n765) );
  XOR2X2 aes_core_keymem_U145 ( .A(aes_core_keymem_n691), .B(
        aes_core_keymem_sboxw[29]), .Y(aes_core_keymem_n757) );
  BUFX12 aes_core_keymem_U144 ( .A(aes_core_keymem_n756), .Y(
        aes_core_keymem_n2407) );
  XOR2X2 aes_core_keymem_U143 ( .A(aes_core_keymem_n733), .B(
        aes_core_keymem_sboxw[8]), .Y(aes_core_keymem_n805) );
  XOR2X2 aes_core_keymem_U142 ( .A(aes_core_keymem_n701), .B(
        aes_core_keymem_sboxw[24]), .Y(aes_core_keymem_n772) );
  BUFX12 aes_core_keymem_U141 ( .A(aes_core_keymem_n771), .Y(
        aes_core_keymem_n2402) );
  XOR2X1 aes_core_keymem_U140 ( .A(aes_core_keymem_prev_key1_reg[126]), .B(
        aes_core_keymem_rcon_reg[6]), .Y(aes_core_keymem_n8) );
  XOR2X1 aes_core_keymem_U139 ( .A(aes_core_keymem_prev_key1_reg[124]), .B(
        aes_core_keymem_rcon_reg[4]), .Y(aes_core_keymem_n7) );
  XOR2X1 aes_core_keymem_U138 ( .A(aes_core_keymem_prev_key1_reg[127]), .B(
        aes_core_keymem_rcon_reg[7]), .Y(aes_core_keymem_n6) );
  XOR2X2 aes_core_keymem_U137 ( .A(aes_core_keymem_n689), .B(
        aes_core_keymem_sboxw[30]), .Y(aes_core_keymem_n754) );
  XOR2X1 aes_core_keymem_U136 ( .A(aes_core_keymem_prev_key1_reg[84]), .B(
        aes_core_keymem_n581), .Y(aes_core_keymem_n645) );
  XOR2X1 aes_core_keymem_U135 ( .A(aes_core_keymem_prev_key1_reg[116]), .B(
        aes_core_new_sboxw[12]), .Y(aes_core_keymem_n581) );
  XOR2X1 aes_core_keymem_U134 ( .A(aes_core_keymem_prev_key1_reg[107]), .B(
        aes_core_new_sboxw[3]), .Y(aes_core_keymem_n599) );
  XOR2X1 aes_core_keymem_U133 ( .A(aes_core_keymem_n731), .B(
        aes_core_keymem_sboxw[9]), .Y(aes_core_keymem_n803) );
  AOI22X1 aes_core_keymem_U132 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n801), .B0(Din[138]), .B1(aes_core_keymem_n2578), .Y(
        aes_core_keymem_n800) );
  XOR2X1 aes_core_keymem_U131 ( .A(aes_core_keymem_n735), .B(
        aes_core_keymem_sboxw[7]), .Y(aes_core_keymem_n807) );
  XOR2X1 aes_core_keymem_U130 ( .A(aes_core_keymem_n699), .B(
        aes_core_keymem_sboxw[25]), .Y(aes_core_keymem_n769) );
  XOR2X1 aes_core_keymem_U129 ( .A(aes_core_keymem_n697), .B(
        aes_core_keymem_sboxw[26]), .Y(aes_core_keymem_n766) );
  BUFX16 aes_core_keymem_U128 ( .A(aes_core_keymem_n765), .Y(
        aes_core_keymem_n2404) );
  XOR2X1 aes_core_keymem_U127 ( .A(aes_core_keymem_prev_key1_reg[95]), .B(
        aes_core_keymem_n558), .Y(aes_core_keymem_n623) );
  XOR2X1 aes_core_keymem_U126 ( .A(aes_core_keymem_prev_key1_reg[92]), .B(
        aes_core_keymem_n565), .Y(aes_core_keymem_n629) );
  XOR2X1 aes_core_keymem_U125 ( .A(aes_core_keymem_prev_key1_reg[91]), .B(
        aes_core_keymem_n567), .Y(aes_core_keymem_n631) );
  XOR2X1 aes_core_keymem_U124 ( .A(aes_core_keymem_prev_key1_reg[87]), .B(
        aes_core_keymem_n575), .Y(aes_core_keymem_n639) );
  XOR2X1 aes_core_keymem_U123 ( .A(aes_core_keymem_prev_key1_reg[86]), .B(
        aes_core_keymem_n577), .Y(aes_core_keymem_n641) );
  XOR2X1 aes_core_keymem_U122 ( .A(aes_core_keymem_prev_key1_reg[83]), .B(
        aes_core_keymem_n583), .Y(aes_core_keymem_n647) );
  XOR2X1 aes_core_keymem_U121 ( .A(aes_core_keymem_prev_key1_reg[82]), .B(
        aes_core_keymem_n585), .Y(aes_core_keymem_n649) );
  XOR2X1 aes_core_keymem_U120 ( .A(aes_core_keymem_prev_key1_reg[81]), .B(
        aes_core_keymem_n587), .Y(aes_core_keymem_n651) );
  XOR2X1 aes_core_keymem_U119 ( .A(aes_core_keymem_prev_key1_reg[80]), .B(
        aes_core_keymem_n589), .Y(aes_core_keymem_n653) );
  XOR2X1 aes_core_keymem_U118 ( .A(aes_core_keymem_prev_key1_reg[79]), .B(
        aes_core_keymem_n591), .Y(aes_core_keymem_n655) );
  XOR2X1 aes_core_keymem_U117 ( .A(aes_core_keymem_prev_key1_reg[76]), .B(
        aes_core_keymem_n597), .Y(aes_core_keymem_n661) );
  XOR2X1 aes_core_keymem_U116 ( .A(aes_core_keymem_prev_key1_reg[75]), .B(
        aes_core_keymem_n599), .Y(aes_core_keymem_n663) );
  XOR2X1 aes_core_keymem_U115 ( .A(aes_core_keymem_prev_key1_reg[74]), .B(
        aes_core_keymem_n601), .Y(aes_core_keymem_n665) );
  XOR2X1 aes_core_keymem_U114 ( .A(aes_core_keymem_prev_key1_reg[119]), .B(
        aes_core_new_sboxw[15]), .Y(aes_core_keymem_n575) );
  XOR2X1 aes_core_keymem_U113 ( .A(aes_core_keymem_prev_key1_reg[115]), .B(
        aes_core_new_sboxw[11]), .Y(aes_core_keymem_n583) );
  XOR2X1 aes_core_keymem_U112 ( .A(aes_core_keymem_prev_key1_reg[114]), .B(
        aes_core_new_sboxw[10]), .Y(aes_core_keymem_n585) );
  XOR2X1 aes_core_keymem_U111 ( .A(aes_core_keymem_prev_key1_reg[113]), .B(
        aes_core_new_sboxw[9]), .Y(aes_core_keymem_n587) );
  XOR2X1 aes_core_keymem_U110 ( .A(aes_core_keymem_prev_key1_reg[112]), .B(
        aes_core_new_sboxw[8]), .Y(aes_core_keymem_n589) );
  XOR2X1 aes_core_keymem_U109 ( .A(aes_core_keymem_prev_key1_reg[111]), .B(
        aes_core_new_sboxw[7]), .Y(aes_core_keymem_n591) );
  XOR2X1 aes_core_keymem_U108 ( .A(aes_core_keymem_prev_key1_reg[108]), .B(
        aes_core_new_sboxw[4]), .Y(aes_core_keymem_n597) );
  XOR2X1 aes_core_keymem_U107 ( .A(aes_core_keymem_prev_key1_reg[106]), .B(
        aes_core_new_sboxw[2]), .Y(aes_core_keymem_n601) );
  XOR2X1 aes_core_keymem_U106 ( .A(aes_core_keymem_prev_key1_reg[100]), .B(
        aes_core_new_sboxw[28]), .Y(aes_core_keymem_n613) );
  XOR2X1 aes_core_keymem_U105 ( .A(aes_core_keymem_prev_key1_reg[103]), .B(
        aes_core_new_sboxw[31]), .Y(aes_core_keymem_n607) );
  XOR2X1 aes_core_keymem_U104 ( .A(aes_core_keymem_prev_key1_reg[99]), .B(
        aes_core_new_sboxw[27]), .Y(aes_core_keymem_n615) );
  XOR2X1 aes_core_keymem_U103 ( .A(aes_core_keymem_prev_key1_reg[97]), .B(
        aes_core_new_sboxw[25]), .Y(aes_core_keymem_n619) );
  XOR2X1 aes_core_keymem_U102 ( .A(aes_core_keymem_prev_key1_reg[118]), .B(
        aes_core_new_sboxw[14]), .Y(aes_core_keymem_n577) );
  BUFX16 aes_core_keymem_U101 ( .A(aes_core_keymem_n818), .Y(
        aes_core_keymem_n544) );
  BUFX16 aes_core_keymem_U100 ( .A(aes_core_keymem_n808), .Y(
        aes_core_keymem_n755) );
  XOR2X1 aes_core_keymem_U99 ( .A(aes_core_keymem_n705), .B(
        aes_core_keymem_sboxw[22]), .Y(aes_core_keymem_n777) );
  XOR2X2 aes_core_keymem_U98 ( .A(aes_core_keymem_prev_key1_reg[96]), .B(
        aes_core_new_sboxw[24]), .Y(aes_core_keymem_n621) );
  XOR2X4 aes_core_keymem_U97 ( .A(aes_core_keymem_prev_key1_reg[69]), .B(
        aes_core_keymem_n611), .Y(aes_core_keymem_n675) );
  XOR2X4 aes_core_keymem_U96 ( .A(aes_core_keymem_prev_key1_reg[70]), .B(
        aes_core_keymem_n609), .Y(aes_core_keymem_n673) );
  XOR2X2 aes_core_keymem_U95 ( .A(aes_core_keymem_prev_key1_reg[68]), .B(
        aes_core_keymem_n613), .Y(aes_core_keymem_n677) );
  XOR2X2 aes_core_keymem_U94 ( .A(aes_core_keymem_prev_key1_reg[71]), .B(
        aes_core_keymem_n607), .Y(aes_core_keymem_n671) );
  XOR2X2 aes_core_keymem_U93 ( .A(aes_core_keymem_prev_key1_reg[67]), .B(
        aes_core_keymem_n615), .Y(aes_core_keymem_n679) );
  XOR2X4 aes_core_keymem_U92 ( .A(aes_core_keymem_prev_key1_reg[64]), .B(
        aes_core_keymem_n621), .Y(aes_core_keymem_n685) );
  INVX1 aes_core_keymem_U91 ( .A(aes_core_keymem_round_ctr_reg[1]), .Y(
        aes_core_keymem_n2768) );
  XOR2X2 aes_core_keymem_U90 ( .A(aes_core_keymem_prev_key1_reg[73]), .B(
        aes_core_keymem_n603), .Y(aes_core_keymem_n667) );
  XOR2X1 aes_core_keymem_U89 ( .A(aes_core_keymem_n15), .B(
        aes_core_new_sboxw[18]), .Y(aes_core_keymem_n569) );
  XOR2X1 aes_core_keymem_U88 ( .A(aes_core_keymem_n11), .B(
        aes_core_new_sboxw[17]), .Y(aes_core_keymem_n571) );
  XOR2X1 aes_core_keymem_U87 ( .A(aes_core_keymem_n8), .B(
        aes_core_new_sboxw[22]), .Y(aes_core_keymem_n561) );
  XOR2X1 aes_core_keymem_U86 ( .A(aes_core_keymem_n10), .B(
        aes_core_new_sboxw[21]), .Y(aes_core_keymem_n563) );
  XOR2X2 aes_core_keymem_U85 ( .A(aes_core_keymem_n713), .B(
        aes_core_keymem_sboxw[18]), .Y(aes_core_keymem_n785) );
  BUFX12 aes_core_keymem_U84 ( .A(aes_core_keymem_n784), .Y(
        aes_core_keymem_n2396) );
  XOR2X2 aes_core_keymem_U83 ( .A(aes_core_keymem_n729), .B(
        aes_core_keymem_sboxw[10]), .Y(aes_core_keymem_n801) );
  BUFX12 aes_core_keymem_U82 ( .A(aes_core_keymem_n798), .Y(
        aes_core_keymem_n770) );
  BUFX12 aes_core_keymem_U81 ( .A(aes_core_keymem_n790), .Y(
        aes_core_keymem_n2393) );
  BUFX12 aes_core_keymem_U80 ( .A(aes_core_keymem_n780), .Y(
        aes_core_keymem_n2398) );
  XOR2X2 aes_core_keymem_U79 ( .A(aes_core_keymem_n7), .B(
        aes_core_new_sboxw[20]), .Y(aes_core_keymem_n565) );
  XOR2X2 aes_core_keymem_U78 ( .A(aes_core_keymem_n6), .B(
        aes_core_new_sboxw[23]), .Y(aes_core_keymem_n558) );
  BUFX8 aes_core_keymem_U77 ( .A(aes_core_keymem_n776), .Y(
        aes_core_keymem_n2400) );
  XOR2X2 aes_core_keymem_U76 ( .A(aes_core_keymem_n687), .B(
        aes_core_keymem_sboxw[31]), .Y(aes_core_keymem_n751) );
  BUFX12 aes_core_keymem_U75 ( .A(aes_core_keymem_n750), .Y(
        aes_core_keymem_n2409) );
  XOR2X2 aes_core_keymem_U74 ( .A(aes_core_keymem_n693), .B(
        aes_core_keymem_sboxw[28]), .Y(aes_core_keymem_n760) );
  BUFX12 aes_core_keymem_U73 ( .A(aes_core_keymem_n759), .Y(
        aes_core_keymem_n2406) );
  XOR2X2 aes_core_keymem_U72 ( .A(aes_core_keymem_prev_key1_reg[89]), .B(
        aes_core_keymem_n571), .Y(aes_core_keymem_n635) );
  XOR2X2 aes_core_keymem_U71 ( .A(aes_core_keymem_prev_key1_reg[90]), .B(
        aes_core_keymem_n569), .Y(aes_core_keymem_n633) );
  XOR2X2 aes_core_keymem_U70 ( .A(aes_core_keymem_prev_key1_reg[94]), .B(
        aes_core_keymem_n561), .Y(aes_core_keymem_n625) );
  XOR2X2 aes_core_keymem_U69 ( .A(aes_core_keymem_prev_key1_reg[93]), .B(
        aes_core_keymem_n563), .Y(aes_core_keymem_n627) );
  XOR2X2 aes_core_keymem_U68 ( .A(aes_core_keymem_n727), .B(
        aes_core_keymem_sboxw[11]), .Y(aes_core_keymem_n799) );
  XOR2X2 aes_core_keymem_U67 ( .A(aes_core_keymem_n715), .B(
        aes_core_keymem_sboxw[17]), .Y(aes_core_keymem_n787) );
  XOR2X2 aes_core_keymem_U66 ( .A(aes_core_keymem_n719), .B(
        aes_core_keymem_sboxw[15]), .Y(aes_core_keymem_n791) );
  XOR2X2 aes_core_keymem_U65 ( .A(aes_core_keymem_n709), .B(
        aes_core_keymem_sboxw[20]), .Y(aes_core_keymem_n781) );
  XOR2X1 aes_core_keymem_U64 ( .A(aes_core_keymem_prev_key1_reg[78]), .B(
        aes_core_keymem_n593), .Y(aes_core_keymem_n657) );
  XOR2X1 aes_core_keymem_U63 ( .A(aes_core_keymem_prev_key1_reg[77]), .B(
        aes_core_keymem_n595), .Y(aes_core_keymem_n659) );
  BUFX16 aes_core_keymem_U62 ( .A(aes_core_keymem_n816), .Y(
        aes_core_keymem_n554) );
  AOI22X4 aes_core_keymem_U61 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n817), .B0(Din[130]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n816) );
  XOR2X1 aes_core_keymem_U60 ( .A(aes_core_keymem_n12), .B(
        aes_core_new_sboxw[16]), .Y(aes_core_keymem_n573) );
  XOR2X1 aes_core_keymem_U59 ( .A(aes_core_keymem_prev_key1_reg[110]), .B(
        aes_core_new_sboxw[6]), .Y(aes_core_keymem_n593) );
  XOR2X1 aes_core_keymem_U58 ( .A(aes_core_keymem_prev_key1_reg[109]), .B(
        aes_core_new_sboxw[5]), .Y(aes_core_keymem_n595) );
  XOR2X2 aes_core_keymem_U57 ( .A(aes_core_keymem_n717), .B(
        aes_core_keymem_sboxw[16]), .Y(aes_core_keymem_n789) );
  XOR2X2 aes_core_keymem_U56 ( .A(aes_core_keymem_prev_key1_reg[88]), .B(
        aes_core_keymem_n573), .Y(aes_core_keymem_n637) );
  XOR2X1 aes_core_keymem_U55 ( .A(aes_core_keymem_prev_key1_reg[104]), .B(
        aes_core_new_sboxw[0]), .Y(aes_core_keymem_n605) );
  XOR2X2 aes_core_keymem_U54 ( .A(aes_core_keymem_prev_key1_reg[72]), .B(
        aes_core_keymem_n605), .Y(aes_core_keymem_n669) );
  OAI221X4 aes_core_keymem_U53 ( .A0(aes_core_keymem_n2765), .A1(
        aes_core_keymem_n821), .B0(aes_core_keymem_key_mem_ctrl_reg[1]), .B1(
        aes_core_keymem_n2773), .C0(aes_core_keymem_n17), .Y(
        aes_core_keymem_n840) );
  DLY1X1 aes_core_keymem_U52 ( .A(aes_core_keymem_n2763), .Y(
        aes_core_keymem_n17) );
  NAND2X1 aes_core_keymem_U51 ( .A(aes_core_enc_round_nr[3]), .B(
        aes_core_enc_round_nr[0]), .Y(aes_core_keymem_n5) );
  NAND2X1 aes_core_keymem_U50 ( .A(aes_core_keymem_n541), .B(
        aes_core_enc_round_nr[3]), .Y(aes_core_keymem_n4) );
  AND3X1 aes_core_keymem_U49 ( .A(aes_core_keymem_n2767), .B(
        aes_core_keymem_n2768), .C(aes_core_keymem_n828), .Y(
        aes_core_keymem_n3) );
  AND3X1 aes_core_keymem_U48 ( .A(aes_core_keymem_n2762), .B(
        aes_core_keymem_n828), .C(aes_core_keymem_n825), .Y(aes_core_keymem_n2) );
  BUFX8 aes_core_keymem_U47 ( .A(aes_core_keymem_n753), .Y(
        aes_core_keymem_n2408) );
  CLKBUFX8 aes_core_keymem_U46 ( .A(aes_core_keymem_n788), .Y(
        aes_core_keymem_n2394) );
  BUFX8 aes_core_keymem_U45 ( .A(aes_core_keymem_n800), .Y(
        aes_core_keymem_n767) );
  BUFX4 aes_core_keymem_U44 ( .A(aes_core_keymem_n804), .Y(
        aes_core_keymem_n761) );
  AOI22X2 aes_core_keymem_U43 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n830), .B0(Din[128]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n820) );
  CLKBUFX8 aes_core_keymem_U42 ( .A(aes_core_keymem_n820), .Y(
        aes_core_keymem_n30) );
  XOR2X1 aes_core_keymem_U41 ( .A(aes_core_keymem_n695), .B(
        aes_core_keymem_sboxw[27]), .Y(aes_core_keymem_n763) );
  CLKBUFX8 aes_core_keymem_U40 ( .A(aes_core_keymem_n762), .Y(
        aes_core_keymem_n2405) );
  BUFX3 aes_core_keymem_U39 ( .A(aes_core_keymem_n768), .Y(
        aes_core_keymem_n2403) );
  XOR2X1 aes_core_keymem_U38 ( .A(aes_core_keymem_n703), .B(
        aes_core_keymem_sboxw[23]), .Y(aes_core_keymem_n775) );
  CLKBUFX8 aes_core_keymem_U37 ( .A(aes_core_keymem_n774), .Y(
        aes_core_keymem_n2401) );
  XOR2X1 aes_core_keymem_U36 ( .A(aes_core_keymem_n707), .B(
        aes_core_keymem_sboxw[21]), .Y(aes_core_keymem_n779) );
  BUFX4 aes_core_keymem_U35 ( .A(aes_core_keymem_n778), .Y(
        aes_core_keymem_n2399) );
  XOR2X1 aes_core_keymem_U34 ( .A(aes_core_keymem_n711), .B(
        aes_core_keymem_sboxw[19]), .Y(aes_core_keymem_n783) );
  CLKBUFX8 aes_core_keymem_U33 ( .A(aes_core_keymem_n782), .Y(
        aes_core_keymem_n2397) );
  CLKBUFX8 aes_core_keymem_U32 ( .A(aes_core_keymem_n786), .Y(
        aes_core_keymem_n2395) );
  XOR2X1 aes_core_keymem_U31 ( .A(aes_core_keymem_n725), .B(
        aes_core_keymem_sboxw[12]), .Y(aes_core_keymem_n797) );
  CLKBUFX8 aes_core_keymem_U30 ( .A(aes_core_keymem_n796), .Y(
        aes_core_keymem_n773) );
  AOI22X1 aes_core_keymem_U29 ( .A0(aes_core_keymem_n2590), .A1(
        aes_core_keymem_n803), .B0(Din[137]), .B1(aes_core_keymem_n2552), .Y(
        aes_core_keymem_n802) );
  BUFX3 aes_core_keymem_U28 ( .A(aes_core_keymem_n802), .Y(
        aes_core_keymem_n764) );
  BUFX4 aes_core_keymem_U27 ( .A(aes_core_keymem_n806), .Y(
        aes_core_keymem_n758) );
  AOI22X2 aes_core_keymem_U26 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n811), .B0(Din[133]), .B1(aes_core_keymem_n2553), .Y(
        aes_core_keymem_n810) );
  BUFX4 aes_core_keymem_U25 ( .A(aes_core_keymem_n810), .Y(
        aes_core_keymem_n752) );
  AOI22X2 aes_core_keymem_U24 ( .A0(aes_core_keymem_n2591), .A1(
        aes_core_keymem_n813), .B0(Din[132]), .B1(aes_core_keymem_n2552), .Y(
        aes_core_keymem_n812) );
  BUFX4 aes_core_keymem_U23 ( .A(aes_core_keymem_n812), .Y(
        aes_core_keymem_n559) );
  XOR2X1 aes_core_keymem_U22 ( .A(aes_core_keymem_n743), .B(
        aes_core_keymem_sboxw[3]), .Y(aes_core_keymem_n815) );
  CLKBUFX8 aes_core_keymem_U21 ( .A(aes_core_keymem_n814), .Y(
        aes_core_keymem_n557) );
  NOR2X1 aes_core_keymem_U20 ( .A(aes_core_keymem_n2767), .B(
        aes_core_keymem_round_ctr_reg[1]), .Y(aes_core_keymem_n824) );
  NOR2X2 aes_core_keymem_U19 ( .A(aes_core_keymem_n2769), .B(
        aes_core_keymem_round_ctr_reg[3]), .Y(aes_core_keymem_n826) );
  NOR2X1 aes_core_keymem_U18 ( .A(aes_core_keymem_n2764), .B(
        aes_core_keymem_round_ctr_reg[2]), .Y(aes_core_keymem_n823) );
  XOR2X1 aes_core_keymem_U17 ( .A(aes_core_keymem_n13), .B(
        aes_core_new_sboxw[19]), .Y(aes_core_keymem_n567) );
  XOR2X1 aes_core_keymem_U16 ( .A(aes_core_keymem_prev_key1_reg[117]), .B(
        aes_core_new_sboxw[13]), .Y(aes_core_keymem_n579) );
  XOR2X1 aes_core_keymem_U15 ( .A(aes_core_keymem_prev_key1_reg[105]), .B(
        aes_core_new_sboxw[1]), .Y(aes_core_keymem_n603) );
  XOR2X2 aes_core_keymem_U14 ( .A(aes_core_keymem_prev_key1_reg[66]), .B(
        aes_core_keymem_n617), .Y(aes_core_keymem_n681) );
  XOR2X1 aes_core_keymem_U13 ( .A(aes_core_keymem_prev_key1_reg[65]), .B(
        aes_core_keymem_n619), .Y(aes_core_keymem_n683) );
  XOR2X2 aes_core_keymem_U12 ( .A(aes_core_keymem_prev_key1_reg[85]), .B(
        aes_core_keymem_n579), .Y(aes_core_keymem_n643) );
  INVX8 aes_core_keymem_U11 ( .A(aes_core_keymem_key_mem_ctrl_reg[0]), .Y(
        aes_core_keymem_n2763) );
  CLKINVX3 aes_core_keymem_U10 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2634) );
  CLKINVX3 aes_core_keymem_U9 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2632) );
  CLKINVX3 aes_core_keymem_U8 ( .A(aes_core_keymem_n2), .Y(
        aes_core_keymem_n2631) );
  CLKINVX3 aes_core_keymem_U7 ( .A(aes_core_keymem_n556), .Y(
        aes_core_keymem_n2608) );
  CLKINVX3 aes_core_keymem_U6 ( .A(aes_core_keymem_n555), .Y(
        aes_core_keymem_n2625) );
  CLKINVX3 aes_core_keymem_U5 ( .A(aes_core_keymem_n829), .Y(
        aes_core_keymem_n2762) );
  CLKINVX3 aes_core_keymem_U4 ( .A(aes_core_keymem_n2556), .Y(
        aes_core_keymem_n2550) );
  NOR2X1 aes_core_keymem_U3 ( .A(aes_core_keymem_n829), .B(
        aes_core_keymem_n2591), .Y(aes_core_keymem_n1) );
  DFFRHQX1 aes_core_keymem_round_ctr_reg_reg_2_ ( .D(aes_core_keymem_n2387), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_round_ctr_reg[2]) );
  DFFRHQX1 aes_core_keymem_round_ctr_reg_reg_3_ ( .D(aes_core_keymem_n2389), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_round_ctr_reg[3]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_0_ ( .D(aes_core_keymem_n2385), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[0]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_2_ ( .D(aes_core_keymem_n2383), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[2]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_5_ ( .D(aes_core_keymem_n2380), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[5]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_6_ ( .D(aes_core_keymem_n2379), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[6]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_3_ ( .D(aes_core_keymem_n2382), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[3]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_7_ ( .D(aes_core_keymem_n2378), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[7]) );
  DFFRHQX1 aes_core_keymem_round_ctr_reg_reg_0_ ( .D(aes_core_keymem_n2386), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_round_ctr_reg[0]) );
  DFFRHQX1 aes_core_keymem_ready_reg_reg ( .D(aes_core_keymem_n841), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_key_ready) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_1_ ( .D(aes_core_keymem_n2384), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[1]) );
  DFFRHQX1 aes_core_keymem_rcon_reg_reg_4_ ( .D(aes_core_keymem_n2381), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_rcon_reg[4]) );
  DFFX4 aes_core_keymem_key_mem_reg_10__126_ ( .D(aes_core_keymem_n854), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[638]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__125_ ( .D(aes_core_keymem_n866), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[637]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__124_ ( .D(aes_core_keymem_n878), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[636]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__123_ ( .D(aes_core_keymem_n890), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[635]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__122_ ( .D(aes_core_keymem_n902), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[634]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__121_ ( .D(aes_core_keymem_n914), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[633]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__120_ ( .D(aes_core_keymem_n926), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[632]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__112_ ( .D(aes_core_keymem_n1022), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[624]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__118_ ( .D(aes_core_keymem_n950), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[630]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__117_ ( .D(aes_core_keymem_n962), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[629]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__116_ ( .D(aes_core_keymem_n974), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[628]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__115_ ( .D(aes_core_keymem_n986), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[627]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__114_ ( .D(aes_core_keymem_n998), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[626]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__113_ ( .D(aes_core_keymem_n1010), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[625]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__108_ ( .D(aes_core_keymem_n1070), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[620]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__111_ ( .D(aes_core_keymem_n1034), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[623]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__110_ ( .D(aes_core_keymem_n1046), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[622]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__109_ ( .D(aes_core_keymem_n1058), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[621]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__106_ ( .D(aes_core_keymem_n1094), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[618]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__107_ ( .D(aes_core_keymem_n1082), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[619]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__105_ ( .D(aes_core_keymem_n1106), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[617]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__104_ ( .D(aes_core_keymem_n1118), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[616]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__103_ ( .D(aes_core_keymem_n1130), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[615]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__96_ ( .D(aes_core_keymem_n1214), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[608]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__102_ ( .D(aes_core_keymem_n1142), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[614]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__101_ ( .D(aes_core_keymem_n1154), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[613]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__100_ ( .D(aes_core_keymem_n1166), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[612]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__99_ ( .D(aes_core_keymem_n1178), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[611]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__98_ ( .D(aes_core_keymem_n1190), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[610]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__97_ ( .D(aes_core_keymem_n1202), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[609]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__87_ ( .D(aes_core_keymem_n1322), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[599]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__95_ ( .D(aes_core_keymem_n1226), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[607]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__94_ ( .D(aes_core_keymem_n1238), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[606]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__93_ ( .D(aes_core_keymem_n1250), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[605]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__92_ ( .D(aes_core_keymem_n1262), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[604]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__91_ ( .D(aes_core_keymem_n1274), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[603]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__90_ ( .D(aes_core_keymem_n1286), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[602]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__89_ ( .D(aes_core_keymem_n1298), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[601]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__88_ ( .D(aes_core_keymem_n1310), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[600]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__80_ ( .D(aes_core_keymem_n1406), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[592]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__86_ ( .D(aes_core_keymem_n1334), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[598]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__85_ ( .D(aes_core_keymem_n1346), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[597]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__84_ ( .D(aes_core_keymem_n1358), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[596]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__83_ ( .D(aes_core_keymem_n1370), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[595]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__82_ ( .D(aes_core_keymem_n1382), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[594]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__81_ ( .D(aes_core_keymem_n1394), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[593]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__76_ ( .D(aes_core_keymem_n1454), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[588]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__79_ ( .D(aes_core_keymem_n1418), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[591]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__78_ ( .D(aes_core_keymem_n1430), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[590]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__77_ ( .D(aes_core_keymem_n1442), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[589]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__74_ ( .D(aes_core_keymem_n1478), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[586]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__75_ ( .D(aes_core_keymem_n1466), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[587]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__73_ ( .D(aes_core_keymem_n1490), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[585]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__72_ ( .D(aes_core_keymem_n1502), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[584]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__71_ ( .D(aes_core_keymem_n1514), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[583]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__64_ ( .D(aes_core_keymem_n1598), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[576]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__70_ ( .D(aes_core_keymem_n1526), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[582]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__69_ ( .D(aes_core_keymem_n1538), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[581]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__68_ ( .D(aes_core_keymem_n1550), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[580]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__67_ ( .D(aes_core_keymem_n1562), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[579]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__66_ ( .D(aes_core_keymem_n1574), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[578]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__65_ ( .D(aes_core_keymem_n1586), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[577]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__55_ ( .D(aes_core_keymem_n1706), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[567]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__63_ ( .D(aes_core_keymem_n1610), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[575]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__62_ ( .D(aes_core_keymem_n1622), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[574]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__61_ ( .D(aes_core_keymem_n1634), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[573]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__60_ ( .D(aes_core_keymem_n1646), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[572]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__59_ ( .D(aes_core_keymem_n1658), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[571]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__58_ ( .D(aes_core_keymem_n1670), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[570]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__57_ ( .D(aes_core_keymem_n1682), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[569]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__56_ ( .D(aes_core_keymem_n1694), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[568]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__48_ ( .D(aes_core_keymem_n1790), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[560]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__54_ ( .D(aes_core_keymem_n1718), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[566]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__53_ ( .D(aes_core_keymem_n1730), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[565]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__52_ ( .D(aes_core_keymem_n1742), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[564]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__51_ ( .D(aes_core_keymem_n1754), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[563]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__50_ ( .D(aes_core_keymem_n1766), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[562]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__49_ ( .D(aes_core_keymem_n1778), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[561]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__44_ ( .D(aes_core_keymem_n1838), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[556]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__47_ ( .D(aes_core_keymem_n1802), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[559]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__46_ ( .D(aes_core_keymem_n1814), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[558]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__45_ ( .D(aes_core_keymem_n1826), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[557]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__42_ ( .D(aes_core_keymem_n1862), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[554]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__43_ ( .D(aes_core_keymem_n1850), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[555]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__41_ ( .D(aes_core_keymem_n1874), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[553]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__40_ ( .D(aes_core_keymem_n1886), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[552]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__39_ ( .D(aes_core_keymem_n1898), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[551]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__32_ ( .D(aes_core_keymem_n1982), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[544]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__38_ ( .D(aes_core_keymem_n1910), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[550]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__37_ ( .D(aes_core_keymem_n1922), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[549]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__36_ ( .D(aes_core_keymem_n1934), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[548]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__35_ ( .D(aes_core_keymem_n1946), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[547]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__34_ ( .D(aes_core_keymem_n1958), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[546]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__33_ ( .D(aes_core_keymem_n1970), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[545]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__23_ ( .D(aes_core_keymem_n2090), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[535]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__31_ ( .D(aes_core_keymem_n1994), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[543]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__30_ ( .D(aes_core_keymem_n2006), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[542]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__29_ ( .D(aes_core_keymem_n2018), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[541]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__28_ ( .D(aes_core_keymem_n2030), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[540]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__27_ ( .D(aes_core_keymem_n2042), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[539]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__26_ ( .D(aes_core_keymem_n2054), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[538]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__25_ ( .D(aes_core_keymem_n2066), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[537]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__24_ ( .D(aes_core_keymem_n2078), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[536]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__16_ ( .D(aes_core_keymem_n2174), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[528]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__22_ ( .D(aes_core_keymem_n2102), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[534]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__21_ ( .D(aes_core_keymem_n2114), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[533]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__20_ ( .D(aes_core_keymem_n2126), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[532]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__19_ ( .D(aes_core_keymem_n2138), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[531]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__18_ ( .D(aes_core_keymem_n2150), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[530]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__17_ ( .D(aes_core_keymem_n2162), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[529]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__12_ ( .D(aes_core_keymem_n2222), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[524]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__15_ ( .D(aes_core_keymem_n2186), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[527]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__14_ ( .D(aes_core_keymem_n2198), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[526]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__13_ ( .D(aes_core_keymem_n2210), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[525]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__10_ ( .D(aes_core_keymem_n2246), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[522]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__11_ ( .D(aes_core_keymem_n2234), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[523]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__9_ ( .D(aes_core_keymem_n2258), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[521]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__8_ ( .D(aes_core_keymem_n2270), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[520]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__7_ ( .D(aes_core_keymem_n2282), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[519]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__0_ ( .D(aes_core_keymem_n2366), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[512]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__6_ ( .D(aes_core_keymem_n2294), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[518]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__5_ ( .D(aes_core_keymem_n2306), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[517]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__4_ ( .D(aes_core_keymem_n2318), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[516]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__3_ ( .D(aes_core_keymem_n2330), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[515]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__2_ ( .D(aes_core_keymem_n2342), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[514]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__1_ ( .D(aes_core_keymem_n2354), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[513]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__119_ ( .D(aes_core_keymem_n938), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[631]), .QN() );
  DFFX4 aes_core_keymem_key_mem_reg_10__127_ ( .D(aes_core_keymem_n842), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[639]), .QN() );
  DFFRHQX1 aes_core_keymem_round_ctr_reg_reg_1_ ( .D(aes_core_keymem_n2761), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_round_ctr_reg[1]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_0_ ( .D(aes_core_keymem_n2377), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[0]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_1_ ( .D(aes_core_keymem_n2365), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[1]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_3_ ( .D(aes_core_keymem_n2341), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[3]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_4_ ( .D(aes_core_keymem_n2329), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[4]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_5_ ( .D(aes_core_keymem_n2317), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[5]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_8_ ( .D(aes_core_keymem_n2281), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[8]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_9_ ( .D(aes_core_keymem_n2269), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[9]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_11_ ( .D(aes_core_keymem_n2245), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[11]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_12_ ( .D(aes_core_keymem_n2233), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[12]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_13_ ( .D(aes_core_keymem_n2221), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[13]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_16_ ( .D(aes_core_keymem_n2185), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[16]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_17_ ( .D(aes_core_keymem_n2173), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[17]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_19_ ( .D(aes_core_keymem_n2149), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[19]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_20_ ( .D(aes_core_keymem_n2137), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[20]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_21_ ( .D(aes_core_keymem_n2125), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[21]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_24_ ( .D(aes_core_keymem_n2089), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[24]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_25_ ( .D(aes_core_keymem_n2077), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[25]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_27_ ( .D(aes_core_keymem_n2053), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[27]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_28_ ( .D(aes_core_keymem_n2041), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[28]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_2_ ( .D(aes_core_keymem_n2353), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[2]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_10_ ( .D(aes_core_keymem_n2257), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[10]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_18_ ( .D(aes_core_keymem_n2161), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[18]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_26_ ( .D(aes_core_keymem_n2065), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[26]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_29_ ( .D(aes_core_keymem_n2029), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[29]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_6_ ( .D(aes_core_keymem_n2305), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[6]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_14_ ( .D(aes_core_keymem_n2209), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[14]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_22_ ( .D(aes_core_keymem_n2113), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[22]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_7_ ( .D(aes_core_keymem_n2293), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[7]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_15_ ( .D(aes_core_keymem_n2197), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[15]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_23_ ( .D(aes_core_keymem_n2101), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[23]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_30_ ( .D(aes_core_keymem_n2017), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[30]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_31_ ( .D(aes_core_keymem_n2005), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_sboxw[31]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__1_ ( .D(aes_core_keymem_n2362), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1025]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__2_ ( .D(aes_core_keymem_n2350), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1026]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__3_ ( .D(aes_core_keymem_n2338), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1027]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__4_ ( .D(aes_core_keymem_n2326), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1028]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__5_ ( .D(aes_core_keymem_n2314), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1029]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__6_ ( .D(aes_core_keymem_n2302), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1030]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__7_ ( .D(aes_core_keymem_n2290), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1031]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__17_ ( .D(aes_core_keymem_n2170), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1041]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__18_ ( .D(aes_core_keymem_n2158), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1042]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__19_ ( .D(aes_core_keymem_n2146), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1043]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__20_ ( .D(aes_core_keymem_n2134), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1044]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__21_ ( .D(aes_core_keymem_n2122), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1045]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__22_ ( .D(aes_core_keymem_n2110), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1046]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__23_ ( .D(aes_core_keymem_n2098), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1047]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__33_ ( .D(aes_core_keymem_n1978), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1057]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__34_ ( .D(aes_core_keymem_n1966), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1058]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__35_ ( .D(aes_core_keymem_n1954), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1059]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__36_ ( .D(aes_core_keymem_n1942), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1060]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__37_ ( .D(aes_core_keymem_n1930), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1061]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__38_ ( .D(aes_core_keymem_n1918), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1062]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__39_ ( .D(aes_core_keymem_n1906), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1063]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__49_ ( .D(aes_core_keymem_n1786), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1073]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__50_ ( .D(aes_core_keymem_n1774), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1074]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__51_ ( .D(aes_core_keymem_n1762), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1075]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__52_ ( .D(aes_core_keymem_n1750), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1076]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__53_ ( .D(aes_core_keymem_n1738), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1077]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__54_ ( .D(aes_core_keymem_n1726), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1078]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__55_ ( .D(aes_core_keymem_n1714), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1079]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__65_ ( .D(aes_core_keymem_n1594), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1089]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__66_ ( .D(aes_core_keymem_n1582), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1090]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__67_ ( .D(aes_core_keymem_n1570), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1091]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__68_ ( .D(aes_core_keymem_n1558), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1092]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__69_ ( .D(aes_core_keymem_n1546), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1093]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__70_ ( .D(aes_core_keymem_n1534), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1094]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__71_ ( .D(aes_core_keymem_n1522), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1095]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__81_ ( .D(aes_core_keymem_n1402), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1105]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__82_ ( .D(aes_core_keymem_n1390), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1106]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__83_ ( .D(aes_core_keymem_n1378), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1107]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__84_ ( .D(aes_core_keymem_n1366), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1108]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__85_ ( .D(aes_core_keymem_n1354), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1109]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__86_ ( .D(aes_core_keymem_n1342), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1110]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__87_ ( .D(aes_core_keymem_n1330), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1111]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__97_ ( .D(aes_core_keymem_n1210), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1121]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__98_ ( .D(aes_core_keymem_n1198), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1122]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__99_ ( .D(aes_core_keymem_n1186), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1123]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__100_ ( .D(aes_core_keymem_n1174), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1124]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__101_ ( .D(aes_core_keymem_n1162), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1125]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__102_ ( .D(aes_core_keymem_n1150), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1126]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__103_ ( .D(aes_core_keymem_n1138), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1127]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__113_ ( .D(aes_core_keymem_n1018), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1137]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__114_ ( .D(aes_core_keymem_n1006), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1138]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__115_ ( .D(aes_core_keymem_n994), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1139]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__116_ ( .D(aes_core_keymem_n982), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1140]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__117_ ( .D(aes_core_keymem_n970), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1141]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__118_ ( .D(aes_core_keymem_n958), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1142]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__119_ ( .D(aes_core_keymem_n946), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1143]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__1_ ( .D(aes_core_keymem_n2361), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[897]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__2_ ( .D(aes_core_keymem_n2349), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[898]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__3_ ( .D(aes_core_keymem_n2337), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[899]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__4_ ( .D(aes_core_keymem_n2325), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[900]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__5_ ( .D(aes_core_keymem_n2313), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[901]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__6_ ( .D(aes_core_keymem_n2301), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[902]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__7_ ( .D(aes_core_keymem_n2289), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[903]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__9_ ( .D(aes_core_keymem_n2265), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[905]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__11_ ( .D(aes_core_keymem_n2241), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[907]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__12_ ( .D(aes_core_keymem_n2229), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[908]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__17_ ( .D(aes_core_keymem_n2169), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[913]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__18_ ( .D(aes_core_keymem_n2157), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[914]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__19_ ( .D(aes_core_keymem_n2145), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[915]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__20_ ( .D(aes_core_keymem_n2133), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[916]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__21_ ( .D(aes_core_keymem_n2121), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[917]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__22_ ( .D(aes_core_keymem_n2109), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[918]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__23_ ( .D(aes_core_keymem_n2097), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[919]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__25_ ( .D(aes_core_keymem_n2073), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[921]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__27_ ( .D(aes_core_keymem_n2049), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[923]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__28_ ( .D(aes_core_keymem_n2037), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[924]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__33_ ( .D(aes_core_keymem_n1977), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[929]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__34_ ( .D(aes_core_keymem_n1965), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[930]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__35_ ( .D(aes_core_keymem_n1953), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[931]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__36_ ( .D(aes_core_keymem_n1941), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[932]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__37_ ( .D(aes_core_keymem_n1929), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[933]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__38_ ( .D(aes_core_keymem_n1917), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[934]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__39_ ( .D(aes_core_keymem_n1905), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[935]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__41_ ( .D(aes_core_keymem_n1881), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[937]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__43_ ( .D(aes_core_keymem_n1857), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[939]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__44_ ( .D(aes_core_keymem_n1845), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[940]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__49_ ( .D(aes_core_keymem_n1785), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[945]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__50_ ( .D(aes_core_keymem_n1773), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[946]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__51_ ( .D(aes_core_keymem_n1761), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[947]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__52_ ( .D(aes_core_keymem_n1749), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[948]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__53_ ( .D(aes_core_keymem_n1737), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[949]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__54_ ( .D(aes_core_keymem_n1725), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[950]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__55_ ( .D(aes_core_keymem_n1713), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[951]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__57_ ( .D(aes_core_keymem_n1689), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[953]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__59_ ( .D(aes_core_keymem_n1665), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[955]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__60_ ( .D(aes_core_keymem_n1653), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[956]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__65_ ( .D(aes_core_keymem_n1593), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[961]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__66_ ( .D(aes_core_keymem_n1581), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[962]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__67_ ( .D(aes_core_keymem_n1569), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[963]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__68_ ( .D(aes_core_keymem_n1557), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[964]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__69_ ( .D(aes_core_keymem_n1545), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[965]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__70_ ( .D(aes_core_keymem_n1533), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[966]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__71_ ( .D(aes_core_keymem_n1521), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[967]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__73_ ( .D(aes_core_keymem_n1497), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[969]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__75_ ( .D(aes_core_keymem_n1473), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[971]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__76_ ( .D(aes_core_keymem_n1461), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[972]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__81_ ( .D(aes_core_keymem_n1401), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[977]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__82_ ( .D(aes_core_keymem_n1389), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[978]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__83_ ( .D(aes_core_keymem_n1377), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[979]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__84_ ( .D(aes_core_keymem_n1365), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[980]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__85_ ( .D(aes_core_keymem_n1353), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[981]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__86_ ( .D(aes_core_keymem_n1341), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[982]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__87_ ( .D(aes_core_keymem_n1329), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[983]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__89_ ( .D(aes_core_keymem_n1305), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[985]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__91_ ( .D(aes_core_keymem_n1281), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[987]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__92_ ( .D(aes_core_keymem_n1269), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[988]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__97_ ( .D(aes_core_keymem_n1209), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[993]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__98_ ( .D(aes_core_keymem_n1197), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[994]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__99_ ( .D(aes_core_keymem_n1185), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[995]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__100_ ( .D(aes_core_keymem_n1173), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[996]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__101_ ( .D(aes_core_keymem_n1161), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[997]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__102_ ( .D(aes_core_keymem_n1149), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[998]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__103_ ( .D(aes_core_keymem_n1137), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[999]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__105_ ( .D(aes_core_keymem_n1113), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1001]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__107_ ( .D(aes_core_keymem_n1089), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1003]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__108_ ( .D(aes_core_keymem_n1077), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1004]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__113_ ( .D(aes_core_keymem_n1017), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1009]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__114_ ( .D(aes_core_keymem_n1005), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1010]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__115_ ( .D(aes_core_keymem_n993), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1011]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__116_ ( .D(aes_core_keymem_n981), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1012]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__117_ ( .D(aes_core_keymem_n969), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1013]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__118_ ( .D(aes_core_keymem_n957), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1014]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__119_ ( .D(aes_core_keymem_n945), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1015]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__121_ ( .D(aes_core_keymem_n921), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1017]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__123_ ( .D(aes_core_keymem_n897), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1019]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__124_ ( .D(aes_core_keymem_n885), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1020]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_120_ ( .D(aes_core_keymem_n937), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[120]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_121_ ( .D(aes_core_keymem_n925), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[121]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_122_ ( .D(aes_core_keymem_n913), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[122]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_123_ ( .D(aes_core_keymem_n901), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[123]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_124_ ( .D(aes_core_keymem_n889), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[124]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_125_ ( .D(aes_core_keymem_n877), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[125]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_126_ ( .D(aes_core_keymem_n865), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[126]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_127_ ( .D(aes_core_keymem_n853), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[127]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__1_ ( .D(aes_core_keymem_n2360), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[385]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__2_ ( .D(aes_core_keymem_n2348), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[386]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__3_ ( .D(aes_core_keymem_n2336), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[387]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__4_ ( .D(aes_core_keymem_n2324), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[388]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__5_ ( .D(aes_core_keymem_n2312), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[389]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__6_ ( .D(aes_core_keymem_n2300), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[390]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__7_ ( .D(aes_core_keymem_n2288), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[391]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__9_ ( .D(aes_core_keymem_n2264), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[393]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__11_ ( .D(aes_core_keymem_n2240), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[395]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__12_ ( .D(aes_core_keymem_n2228), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[396]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__17_ ( .D(aes_core_keymem_n2168), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[401]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__18_ ( .D(aes_core_keymem_n2156), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[402]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__19_ ( .D(aes_core_keymem_n2144), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[403]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__20_ ( .D(aes_core_keymem_n2132), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[404]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__21_ ( .D(aes_core_keymem_n2120), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[405]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__22_ ( .D(aes_core_keymem_n2108), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[406]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__23_ ( .D(aes_core_keymem_n2096), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[407]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__33_ ( .D(aes_core_keymem_n1976), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[417]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__34_ ( .D(aes_core_keymem_n1964), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[418]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__35_ ( .D(aes_core_keymem_n1952), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[419]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__36_ ( .D(aes_core_keymem_n1940), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[420]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__37_ ( .D(aes_core_keymem_n1928), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[421]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__38_ ( .D(aes_core_keymem_n1916), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[422]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__39_ ( .D(aes_core_keymem_n1904), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[423]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__41_ ( .D(aes_core_keymem_n1880), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[425]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__43_ ( .D(aes_core_keymem_n1856), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[427]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__44_ ( .D(aes_core_keymem_n1844), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[428]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__49_ ( .D(aes_core_keymem_n1784), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[433]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__50_ ( .D(aes_core_keymem_n1772), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[434]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__51_ ( .D(aes_core_keymem_n1760), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[435]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__52_ ( .D(aes_core_keymem_n1748), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[436]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__53_ ( .D(aes_core_keymem_n1736), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[437]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__54_ ( .D(aes_core_keymem_n1724), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[438]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__55_ ( .D(aes_core_keymem_n1712), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[439]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__65_ ( .D(aes_core_keymem_n1592), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[449]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__66_ ( .D(aes_core_keymem_n1580), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[450]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__67_ ( .D(aes_core_keymem_n1568), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[451]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__68_ ( .D(aes_core_keymem_n1556), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[452]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__69_ ( .D(aes_core_keymem_n1544), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[453]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__70_ ( .D(aes_core_keymem_n1532), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[454]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__71_ ( .D(aes_core_keymem_n1520), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[455]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__73_ ( .D(aes_core_keymem_n1496), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[457]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__75_ ( .D(aes_core_keymem_n1472), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[459]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__76_ ( .D(aes_core_keymem_n1460), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[460]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__81_ ( .D(aes_core_keymem_n1400), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[465]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__82_ ( .D(aes_core_keymem_n1388), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[466]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__83_ ( .D(aes_core_keymem_n1376), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[467]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__84_ ( .D(aes_core_keymem_n1364), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[468]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__85_ ( .D(aes_core_keymem_n1352), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[469]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__86_ ( .D(aes_core_keymem_n1340), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[470]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__87_ ( .D(aes_core_keymem_n1328), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[471]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__97_ ( .D(aes_core_keymem_n1208), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[481]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__98_ ( .D(aes_core_keymem_n1196), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[482]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__99_ ( .D(aes_core_keymem_n1184), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[483]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__100_ ( .D(aes_core_keymem_n1172), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[484]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__101_ ( .D(aes_core_keymem_n1160), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[485]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__102_ ( .D(aes_core_keymem_n1148), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[486]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__103_ ( .D(aes_core_keymem_n1136), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[487]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__105_ ( .D(aes_core_keymem_n1112), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[489]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__107_ ( .D(aes_core_keymem_n1088), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[491]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__108_ ( .D(aes_core_keymem_n1076), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[492]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__113_ ( .D(aes_core_keymem_n1016), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[497]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__114_ ( .D(aes_core_keymem_n1004), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[498]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__115_ ( .D(aes_core_keymem_n992), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[499]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__116_ ( .D(aes_core_keymem_n980), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[500]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__117_ ( .D(aes_core_keymem_n968), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[501]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__118_ ( .D(aes_core_keymem_n956), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[502]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__119_ ( .D(aes_core_keymem_n944), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[503]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__1_ ( .D(aes_core_keymem_n2357), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[1]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__2_ ( .D(aes_core_keymem_n2345), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[2]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__3_ ( .D(aes_core_keymem_n2333), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[3]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__4_ ( .D(aes_core_keymem_n2321), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[4]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__5_ ( .D(aes_core_keymem_n2309), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[5]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__6_ ( .D(aes_core_keymem_n2297), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[6]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__7_ ( .D(aes_core_keymem_n2285), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[7]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__9_ ( .D(aes_core_keymem_n2261), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[9]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__11_ ( .D(aes_core_keymem_n2237), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[11]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__12_ ( .D(aes_core_keymem_n2225), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[12]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__17_ ( .D(aes_core_keymem_n2165), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[17]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__18_ ( .D(aes_core_keymem_n2153), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[18]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__19_ ( .D(aes_core_keymem_n2141), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[19]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__20_ ( .D(aes_core_keymem_n2129), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[20]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__21_ ( .D(aes_core_keymem_n2117), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[21]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__22_ ( .D(aes_core_keymem_n2105), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[22]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__23_ ( .D(aes_core_keymem_n2093), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[23]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__33_ ( .D(aes_core_keymem_n1973), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[33]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__34_ ( .D(aes_core_keymem_n1961), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[34]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__35_ ( .D(aes_core_keymem_n1949), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[35]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__36_ ( .D(aes_core_keymem_n1937), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[36]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__37_ ( .D(aes_core_keymem_n1925), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[37]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__38_ ( .D(aes_core_keymem_n1913), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[38]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__39_ ( .D(aes_core_keymem_n1901), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[39]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__41_ ( .D(aes_core_keymem_n1877), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[41]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__43_ ( .D(aes_core_keymem_n1853), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[43]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__44_ ( .D(aes_core_keymem_n1841), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[44]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__49_ ( .D(aes_core_keymem_n1781), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[49]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__50_ ( .D(aes_core_keymem_n1769), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[50]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__51_ ( .D(aes_core_keymem_n1757), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[51]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__52_ ( .D(aes_core_keymem_n1745), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[52]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__53_ ( .D(aes_core_keymem_n1733), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[53]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__54_ ( .D(aes_core_keymem_n1721), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[54]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__55_ ( .D(aes_core_keymem_n1709), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[55]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__65_ ( .D(aes_core_keymem_n1589), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[65]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__66_ ( .D(aes_core_keymem_n1577), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[66]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__67_ ( .D(aes_core_keymem_n1565), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[67]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__68_ ( .D(aes_core_keymem_n1553), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[68]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__69_ ( .D(aes_core_keymem_n1541), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[69]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__70_ ( .D(aes_core_keymem_n1529), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[70]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__71_ ( .D(aes_core_keymem_n1517), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[71]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__73_ ( .D(aes_core_keymem_n1493), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[73]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__75_ ( .D(aes_core_keymem_n1469), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[75]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__76_ ( .D(aes_core_keymem_n1457), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[76]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__81_ ( .D(aes_core_keymem_n1397), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[81]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__82_ ( .D(aes_core_keymem_n1385), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[82]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__83_ ( .D(aes_core_keymem_n1373), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[83]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__84_ ( .D(aes_core_keymem_n1361), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[84]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__85_ ( .D(aes_core_keymem_n1349), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[85]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__86_ ( .D(aes_core_keymem_n1337), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[86]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__87_ ( .D(aes_core_keymem_n1325), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[87]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__97_ ( .D(aes_core_keymem_n1205), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[97]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__98_ ( .D(aes_core_keymem_n1193), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[98]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__99_ ( .D(aes_core_keymem_n1181), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[99]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__100_ ( .D(aes_core_keymem_n1169), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[100]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__101_ ( .D(aes_core_keymem_n1157), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[101]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__102_ ( .D(aes_core_keymem_n1145), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[102]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__103_ ( .D(aes_core_keymem_n1133), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[103]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__105_ ( .D(aes_core_keymem_n1109), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[105]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__107_ ( .D(aes_core_keymem_n1085), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[107]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__108_ ( .D(aes_core_keymem_n1073), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[108]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__113_ ( .D(aes_core_keymem_n1013), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[113]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__114_ ( .D(aes_core_keymem_n1001), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[114]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__115_ ( .D(aes_core_keymem_n989), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[115]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__116_ ( .D(aes_core_keymem_n977), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[116]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__117_ ( .D(aes_core_keymem_n965), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[117]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__118_ ( .D(aes_core_keymem_n953), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[118]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__119_ ( .D(aes_core_keymem_n941), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[119]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__1_ ( .D(aes_core_keymem_n2358), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[129]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__2_ ( .D(aes_core_keymem_n2346), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[130]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__3_ ( .D(aes_core_keymem_n2334), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[131]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__4_ ( .D(aes_core_keymem_n2322), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[132]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__5_ ( .D(aes_core_keymem_n2310), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[133]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__6_ ( .D(aes_core_keymem_n2298), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[134]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__7_ ( .D(aes_core_keymem_n2286), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[135]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__9_ ( .D(aes_core_keymem_n2262), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[137]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__11_ ( .D(aes_core_keymem_n2238), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[139]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__12_ ( .D(aes_core_keymem_n2226), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[140]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__17_ ( .D(aes_core_keymem_n2166), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[145]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__18_ ( .D(aes_core_keymem_n2154), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[146]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__19_ ( .D(aes_core_keymem_n2142), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[147]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__20_ ( .D(aes_core_keymem_n2130), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[148]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__21_ ( .D(aes_core_keymem_n2118), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[149]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__22_ ( .D(aes_core_keymem_n2106), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[150]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__23_ ( .D(aes_core_keymem_n2094), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[151]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__25_ ( .D(aes_core_keymem_n2070), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[153]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__27_ ( .D(aes_core_keymem_n2046), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[155]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__28_ ( .D(aes_core_keymem_n2034), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[156]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__33_ ( .D(aes_core_keymem_n1974), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[161]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__34_ ( .D(aes_core_keymem_n1962), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[162]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__35_ ( .D(aes_core_keymem_n1950), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[163]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__36_ ( .D(aes_core_keymem_n1938), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[164]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__37_ ( .D(aes_core_keymem_n1926), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[165]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__38_ ( .D(aes_core_keymem_n1914), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[166]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__39_ ( .D(aes_core_keymem_n1902), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[167]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__41_ ( .D(aes_core_keymem_n1878), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[169]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__43_ ( .D(aes_core_keymem_n1854), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[171]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__44_ ( .D(aes_core_keymem_n1842), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[172]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__49_ ( .D(aes_core_keymem_n1782), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[177]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__50_ ( .D(aes_core_keymem_n1770), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[178]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__51_ ( .D(aes_core_keymem_n1758), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[179]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__52_ ( .D(aes_core_keymem_n1746), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[180]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__53_ ( .D(aes_core_keymem_n1734), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[181]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__54_ ( .D(aes_core_keymem_n1722), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[182]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__55_ ( .D(aes_core_keymem_n1710), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[183]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__57_ ( .D(aes_core_keymem_n1686), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[185]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__59_ ( .D(aes_core_keymem_n1662), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[187]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__60_ ( .D(aes_core_keymem_n1650), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[188]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__65_ ( .D(aes_core_keymem_n1590), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[193]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__66_ ( .D(aes_core_keymem_n1578), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[194]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__67_ ( .D(aes_core_keymem_n1566), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[195]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__68_ ( .D(aes_core_keymem_n1554), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[196]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__69_ ( .D(aes_core_keymem_n1542), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[197]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__70_ ( .D(aes_core_keymem_n1530), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[198]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__71_ ( .D(aes_core_keymem_n1518), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[199]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__73_ ( .D(aes_core_keymem_n1494), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[201]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__75_ ( .D(aes_core_keymem_n1470), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[203]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__76_ ( .D(aes_core_keymem_n1458), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[204]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__81_ ( .D(aes_core_keymem_n1398), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[209]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__82_ ( .D(aes_core_keymem_n1386), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[210]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__83_ ( .D(aes_core_keymem_n1374), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[211]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__84_ ( .D(aes_core_keymem_n1362), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[212]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__85_ ( .D(aes_core_keymem_n1350), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[213]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__86_ ( .D(aes_core_keymem_n1338), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[214]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__87_ ( .D(aes_core_keymem_n1326), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[215]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__89_ ( .D(aes_core_keymem_n1302), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[217]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__91_ ( .D(aes_core_keymem_n1278), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[219]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__92_ ( .D(aes_core_keymem_n1266), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[220]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__97_ ( .D(aes_core_keymem_n1206), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[225]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__98_ ( .D(aes_core_keymem_n1194), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[226]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__99_ ( .D(aes_core_keymem_n1182), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[227]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__100_ ( .D(aes_core_keymem_n1170), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[228]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__101_ ( .D(aes_core_keymem_n1158), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[229]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__102_ ( .D(aes_core_keymem_n1146), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[230]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__103_ ( .D(aes_core_keymem_n1134), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[231]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__105_ ( .D(aes_core_keymem_n1110), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[233]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__107_ ( .D(aes_core_keymem_n1086), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[235]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__108_ ( .D(aes_core_keymem_n1074), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[236]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__113_ ( .D(aes_core_keymem_n1014), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[241]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__114_ ( .D(aes_core_keymem_n1002), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[242]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__115_ ( .D(aes_core_keymem_n990), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[243]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__116_ ( .D(aes_core_keymem_n978), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[244]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__117_ ( .D(aes_core_keymem_n966), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[245]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__118_ ( .D(aes_core_keymem_n954), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[246]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__119_ ( .D(aes_core_keymem_n942), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[247]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__121_ ( .D(aes_core_keymem_n918), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[249]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__123_ ( .D(aes_core_keymem_n894), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[251]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__124_ ( .D(aes_core_keymem_n882), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[252]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__1_ ( .D(aes_core_keymem_n2355), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[641]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__2_ ( .D(aes_core_keymem_n2343), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[642]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__3_ ( .D(aes_core_keymem_n2331), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[643]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__4_ ( .D(aes_core_keymem_n2319), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[644]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__5_ ( .D(aes_core_keymem_n2307), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[645]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__6_ ( .D(aes_core_keymem_n2295), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[646]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__7_ ( .D(aes_core_keymem_n2283), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[647]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__9_ ( .D(aes_core_keymem_n2259), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[649]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__11_ ( .D(aes_core_keymem_n2235), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[651]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__12_ ( .D(aes_core_keymem_n2223), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[652]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__17_ ( .D(aes_core_keymem_n2163), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[657]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__18_ ( .D(aes_core_keymem_n2151), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[658]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__19_ ( .D(aes_core_keymem_n2139), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[659]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__20_ ( .D(aes_core_keymem_n2127), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[660]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__21_ ( .D(aes_core_keymem_n2115), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[661]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__22_ ( .D(aes_core_keymem_n2103), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[662]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__23_ ( .D(aes_core_keymem_n2091), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[663]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__25_ ( .D(aes_core_keymem_n2067), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[665]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__27_ ( .D(aes_core_keymem_n2043), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[667]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__28_ ( .D(aes_core_keymem_n2031), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[668]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__33_ ( .D(aes_core_keymem_n1971), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[673]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__34_ ( .D(aes_core_keymem_n1959), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[674]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__35_ ( .D(aes_core_keymem_n1947), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[675]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__36_ ( .D(aes_core_keymem_n1935), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[676]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__37_ ( .D(aes_core_keymem_n1923), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[677]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__38_ ( .D(aes_core_keymem_n1911), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[678]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__39_ ( .D(aes_core_keymem_n1899), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[679]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__41_ ( .D(aes_core_keymem_n1875), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[681]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__43_ ( .D(aes_core_keymem_n1851), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[683]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__44_ ( .D(aes_core_keymem_n1839), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[684]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__49_ ( .D(aes_core_keymem_n1779), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[689]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__50_ ( .D(aes_core_keymem_n1767), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[690]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__51_ ( .D(aes_core_keymem_n1755), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[691]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__52_ ( .D(aes_core_keymem_n1743), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[692]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__53_ ( .D(aes_core_keymem_n1731), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[693]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__54_ ( .D(aes_core_keymem_n1719), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[694]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__55_ ( .D(aes_core_keymem_n1707), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[695]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__57_ ( .D(aes_core_keymem_n1683), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[697]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__59_ ( .D(aes_core_keymem_n1659), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[699]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__60_ ( .D(aes_core_keymem_n1647), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[700]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__65_ ( .D(aes_core_keymem_n1587), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[705]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__66_ ( .D(aes_core_keymem_n1575), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[706]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__67_ ( .D(aes_core_keymem_n1563), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[707]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__68_ ( .D(aes_core_keymem_n1551), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[708]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__69_ ( .D(aes_core_keymem_n1539), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[709]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__70_ ( .D(aes_core_keymem_n1527), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[710]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__71_ ( .D(aes_core_keymem_n1515), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[711]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__73_ ( .D(aes_core_keymem_n1491), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[713]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__75_ ( .D(aes_core_keymem_n1467), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[715]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__76_ ( .D(aes_core_keymem_n1455), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[716]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__81_ ( .D(aes_core_keymem_n1395), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[721]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__82_ ( .D(aes_core_keymem_n1383), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[722]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__83_ ( .D(aes_core_keymem_n1371), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[723]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__84_ ( .D(aes_core_keymem_n1359), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[724]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__85_ ( .D(aes_core_keymem_n1347), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[725]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__86_ ( .D(aes_core_keymem_n1335), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[726]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__87_ ( .D(aes_core_keymem_n1323), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[727]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__89_ ( .D(aes_core_keymem_n1299), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[729]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__91_ ( .D(aes_core_keymem_n1275), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[731]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__92_ ( .D(aes_core_keymem_n1263), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[732]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__97_ ( .D(aes_core_keymem_n1203), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[737]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__98_ ( .D(aes_core_keymem_n1191), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[738]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__99_ ( .D(aes_core_keymem_n1179), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[739]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__100_ ( .D(aes_core_keymem_n1167), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[740]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__101_ ( .D(aes_core_keymem_n1155), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[741]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__102_ ( .D(aes_core_keymem_n1143), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[742]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__103_ ( .D(aes_core_keymem_n1131), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[743]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__105_ ( .D(aes_core_keymem_n1107), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[745]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__107_ ( .D(aes_core_keymem_n1083), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[747]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__108_ ( .D(aes_core_keymem_n1071), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[748]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__113_ ( .D(aes_core_keymem_n1011), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[753]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__114_ ( .D(aes_core_keymem_n999), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[754]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__115_ ( .D(aes_core_keymem_n987), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[755]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__116_ ( .D(aes_core_keymem_n975), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[756]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__117_ ( .D(aes_core_keymem_n963), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[757]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__118_ ( .D(aes_core_keymem_n951), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[758]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__119_ ( .D(aes_core_keymem_n939), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[759]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__121_ ( .D(aes_core_keymem_n915), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[761]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__123_ ( .D(aes_core_keymem_n891), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[763]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__124_ ( .D(aes_core_keymem_n879), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[764]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__0_ ( .D(aes_core_keymem_n2375), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1152]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__1_ ( .D(aes_core_keymem_n2363), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1153]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__2_ ( .D(aes_core_keymem_n2351), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1154]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__3_ ( .D(aes_core_keymem_n2339), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1155]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__4_ ( .D(aes_core_keymem_n2327), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1156]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__5_ ( .D(aes_core_keymem_n2315), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1157]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__6_ ( .D(aes_core_keymem_n2303), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1158]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__7_ ( .D(aes_core_keymem_n2291), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1159]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__8_ ( .D(aes_core_keymem_n2279), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1160]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__9_ ( .D(aes_core_keymem_n2267), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1161]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__10_ ( .D(aes_core_keymem_n2255), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1162]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__11_ ( .D(aes_core_keymem_n2243), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1163]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__12_ ( .D(aes_core_keymem_n2231), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1164]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__13_ ( .D(aes_core_keymem_n2219), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1165]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__14_ ( .D(aes_core_keymem_n2207), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1166]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__15_ ( .D(aes_core_keymem_n2195), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1167]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__16_ ( .D(aes_core_keymem_n2183), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1168]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__17_ ( .D(aes_core_keymem_n2171), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1169]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__18_ ( .D(aes_core_keymem_n2159), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1170]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__19_ ( .D(aes_core_keymem_n2147), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1171]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__20_ ( .D(aes_core_keymem_n2135), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1172]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__21_ ( .D(aes_core_keymem_n2123), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1173]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__22_ ( .D(aes_core_keymem_n2111), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1174]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__23_ ( .D(aes_core_keymem_n2099), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1175]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__24_ ( .D(aes_core_keymem_n2087), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1176]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__25_ ( .D(aes_core_keymem_n2075), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1177]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__26_ ( .D(aes_core_keymem_n2063), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1178]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__27_ ( .D(aes_core_keymem_n2051), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1179]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__28_ ( .D(aes_core_keymem_n2039), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1180]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__29_ ( .D(aes_core_keymem_n2027), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1181]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__30_ ( .D(aes_core_keymem_n2015), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1182]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__31_ ( .D(aes_core_keymem_n2003), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1183]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__32_ ( .D(aes_core_keymem_n1991), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1184]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__33_ ( .D(aes_core_keymem_n1979), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1185]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__34_ ( .D(aes_core_keymem_n1967), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1186]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__35_ ( .D(aes_core_keymem_n1955), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1187]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__36_ ( .D(aes_core_keymem_n1943), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1188]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__37_ ( .D(aes_core_keymem_n1931), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1189]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__38_ ( .D(aes_core_keymem_n1919), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1190]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__39_ ( .D(aes_core_keymem_n1907), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1191]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__40_ ( .D(aes_core_keymem_n1895), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1192]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__41_ ( .D(aes_core_keymem_n1883), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1193]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__42_ ( .D(aes_core_keymem_n1871), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1194]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__43_ ( .D(aes_core_keymem_n1859), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1195]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__44_ ( .D(aes_core_keymem_n1847), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1196]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__45_ ( .D(aes_core_keymem_n1835), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1197]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__46_ ( .D(aes_core_keymem_n1823), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1198]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__47_ ( .D(aes_core_keymem_n1811), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1199]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__48_ ( .D(aes_core_keymem_n1799), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1200]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__49_ ( .D(aes_core_keymem_n1787), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1201]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__50_ ( .D(aes_core_keymem_n1775), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1202]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__51_ ( .D(aes_core_keymem_n1763), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1203]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__52_ ( .D(aes_core_keymem_n1751), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1204]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__53_ ( .D(aes_core_keymem_n1739), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1205]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__54_ ( .D(aes_core_keymem_n1727), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1206]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__55_ ( .D(aes_core_keymem_n1715), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1207]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__56_ ( .D(aes_core_keymem_n1703), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1208]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__57_ ( .D(aes_core_keymem_n1691), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1209]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__58_ ( .D(aes_core_keymem_n1679), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1210]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__59_ ( .D(aes_core_keymem_n1667), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1211]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__60_ ( .D(aes_core_keymem_n1655), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1212]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__61_ ( .D(aes_core_keymem_n1643), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1213]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__62_ ( .D(aes_core_keymem_n1631), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1214]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__63_ ( .D(aes_core_keymem_n1619), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1215]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__64_ ( .D(aes_core_keymem_n1607), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1216]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__65_ ( .D(aes_core_keymem_n1595), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1217]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__66_ ( .D(aes_core_keymem_n1583), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1218]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__67_ ( .D(aes_core_keymem_n1571), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1219]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__68_ ( .D(aes_core_keymem_n1559), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1220]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__69_ ( .D(aes_core_keymem_n1547), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1221]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__70_ ( .D(aes_core_keymem_n1535), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1222]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__71_ ( .D(aes_core_keymem_n1523), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1223]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__72_ ( .D(aes_core_keymem_n1511), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1224]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__73_ ( .D(aes_core_keymem_n1499), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1225]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__74_ ( .D(aes_core_keymem_n1487), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1226]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__75_ ( .D(aes_core_keymem_n1475), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1227]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__76_ ( .D(aes_core_keymem_n1463), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1228]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__77_ ( .D(aes_core_keymem_n1451), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1229]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__78_ ( .D(aes_core_keymem_n1439), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1230]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__79_ ( .D(aes_core_keymem_n1427), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1231]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__80_ ( .D(aes_core_keymem_n1415), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1232]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__81_ ( .D(aes_core_keymem_n1403), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1233]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__82_ ( .D(aes_core_keymem_n1391), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1234]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__83_ ( .D(aes_core_keymem_n1379), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1235]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__84_ ( .D(aes_core_keymem_n1367), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1236]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__85_ ( .D(aes_core_keymem_n1355), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1237]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__86_ ( .D(aes_core_keymem_n1343), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1238]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__87_ ( .D(aes_core_keymem_n1331), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1239]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__88_ ( .D(aes_core_keymem_n1319), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1240]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__89_ ( .D(aes_core_keymem_n1307), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1241]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__90_ ( .D(aes_core_keymem_n1295), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1242]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__91_ ( .D(aes_core_keymem_n1283), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1243]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__92_ ( .D(aes_core_keymem_n1271), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1244]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__93_ ( .D(aes_core_keymem_n1259), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1245]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__94_ ( .D(aes_core_keymem_n1247), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1246]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__95_ ( .D(aes_core_keymem_n1235), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1247]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__96_ ( .D(aes_core_keymem_n1223), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1248]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__97_ ( .D(aes_core_keymem_n1211), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1249]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__98_ ( .D(aes_core_keymem_n1199), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1250]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__99_ ( .D(aes_core_keymem_n1187), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1251]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__100_ ( .D(aes_core_keymem_n1175), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1252]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__101_ ( .D(aes_core_keymem_n1163), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1253]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__102_ ( .D(aes_core_keymem_n1151), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1254]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__103_ ( .D(aes_core_keymem_n1139), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1255]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__104_ ( .D(aes_core_keymem_n1127), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1256]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__105_ ( .D(aes_core_keymem_n1115), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1257]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__106_ ( .D(aes_core_keymem_n1103), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1258]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__107_ ( .D(aes_core_keymem_n1091), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1259]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__108_ ( .D(aes_core_keymem_n1079), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1260]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__109_ ( .D(aes_core_keymem_n1067), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1261]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__110_ ( .D(aes_core_keymem_n1055), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1262]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__111_ ( .D(aes_core_keymem_n1043), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1263]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__112_ ( .D(aes_core_keymem_n1031), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1264]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__113_ ( .D(aes_core_keymem_n1019), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1265]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__114_ ( .D(aes_core_keymem_n1007), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1266]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__115_ ( .D(aes_core_keymem_n995), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1267]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__116_ ( .D(aes_core_keymem_n983), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1268]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__117_ ( .D(aes_core_keymem_n971), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1269]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__118_ ( .D(aes_core_keymem_n959), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1270]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__119_ ( .D(aes_core_keymem_n947), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1271]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__120_ ( .D(aes_core_keymem_n935), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1272]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__121_ ( .D(aes_core_keymem_n923), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1273]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__122_ ( .D(aes_core_keymem_n911), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1274]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__123_ ( .D(aes_core_keymem_n899), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1275]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__124_ ( .D(aes_core_keymem_n887), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1276]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__125_ ( .D(aes_core_keymem_n875), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1277]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__126_ ( .D(aes_core_keymem_n863), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1278]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_1__127_ ( .D(aes_core_keymem_n851), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1279]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__0_ ( .D(aes_core_keymem_n2376), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1280]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__1_ ( .D(aes_core_keymem_n2364), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1281]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__2_ ( .D(aes_core_keymem_n2352), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1282]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__3_ ( .D(aes_core_keymem_n2340), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1283]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__4_ ( .D(aes_core_keymem_n2328), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1284]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__5_ ( .D(aes_core_keymem_n2316), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1285]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__6_ ( .D(aes_core_keymem_n2304), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1286]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__7_ ( .D(aes_core_keymem_n2292), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1287]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__8_ ( .D(aes_core_keymem_n2280), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1288]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__9_ ( .D(aes_core_keymem_n2268), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1289]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__10_ ( .D(aes_core_keymem_n2256), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1290]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__11_ ( .D(aes_core_keymem_n2244), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1291]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__12_ ( .D(aes_core_keymem_n2232), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1292]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__13_ ( .D(aes_core_keymem_n2220), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1293]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__14_ ( .D(aes_core_keymem_n2208), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1294]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__15_ ( .D(aes_core_keymem_n2196), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1295]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__16_ ( .D(aes_core_keymem_n2184), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1296]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__17_ ( .D(aes_core_keymem_n2172), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1297]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__18_ ( .D(aes_core_keymem_n2160), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1298]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__19_ ( .D(aes_core_keymem_n2148), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1299]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__20_ ( .D(aes_core_keymem_n2136), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1300]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__21_ ( .D(aes_core_keymem_n2124), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1301]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__22_ ( .D(aes_core_keymem_n2112), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1302]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__23_ ( .D(aes_core_keymem_n2100), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1303]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__24_ ( .D(aes_core_keymem_n2088), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1304]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__25_ ( .D(aes_core_keymem_n2076), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1305]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__26_ ( .D(aes_core_keymem_n2064), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1306]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__27_ ( .D(aes_core_keymem_n2052), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1307]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__28_ ( .D(aes_core_keymem_n2040), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1308]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__29_ ( .D(aes_core_keymem_n2028), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1309]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__30_ ( .D(aes_core_keymem_n2016), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1310]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__31_ ( .D(aes_core_keymem_n2004), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1311]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__32_ ( .D(aes_core_keymem_n1992), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1312]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__33_ ( .D(aes_core_keymem_n1980), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1313]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__34_ ( .D(aes_core_keymem_n1968), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1314]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__35_ ( .D(aes_core_keymem_n1956), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1315]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__36_ ( .D(aes_core_keymem_n1944), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1316]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__37_ ( .D(aes_core_keymem_n1932), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1317]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__38_ ( .D(aes_core_keymem_n1920), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1318]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__39_ ( .D(aes_core_keymem_n1908), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1319]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__40_ ( .D(aes_core_keymem_n1896), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1320]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__41_ ( .D(aes_core_keymem_n1884), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1321]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__42_ ( .D(aes_core_keymem_n1872), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1322]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__43_ ( .D(aes_core_keymem_n1860), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1323]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__44_ ( .D(aes_core_keymem_n1848), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1324]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__45_ ( .D(aes_core_keymem_n1836), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1325]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__46_ ( .D(aes_core_keymem_n1824), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1326]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__47_ ( .D(aes_core_keymem_n1812), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1327]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__48_ ( .D(aes_core_keymem_n1800), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1328]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__49_ ( .D(aes_core_keymem_n1788), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1329]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__50_ ( .D(aes_core_keymem_n1776), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1330]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__51_ ( .D(aes_core_keymem_n1764), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1331]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__52_ ( .D(aes_core_keymem_n1752), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1332]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__53_ ( .D(aes_core_keymem_n1740), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1333]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__54_ ( .D(aes_core_keymem_n1728), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1334]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__55_ ( .D(aes_core_keymem_n1716), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1335]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__56_ ( .D(aes_core_keymem_n1704), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1336]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__57_ ( .D(aes_core_keymem_n1692), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1337]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__58_ ( .D(aes_core_keymem_n1680), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1338]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__59_ ( .D(aes_core_keymem_n1668), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1339]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__60_ ( .D(aes_core_keymem_n1656), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1340]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__61_ ( .D(aes_core_keymem_n1644), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1341]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__62_ ( .D(aes_core_keymem_n1632), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1342]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__63_ ( .D(aes_core_keymem_n1620), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1343]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__64_ ( .D(aes_core_keymem_n1608), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1344]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__65_ ( .D(aes_core_keymem_n1596), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1345]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__66_ ( .D(aes_core_keymem_n1584), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1346]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__67_ ( .D(aes_core_keymem_n1572), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1347]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__68_ ( .D(aes_core_keymem_n1560), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1348]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__69_ ( .D(aes_core_keymem_n1548), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1349]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__70_ ( .D(aes_core_keymem_n1536), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1350]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__71_ ( .D(aes_core_keymem_n1524), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1351]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__72_ ( .D(aes_core_keymem_n1512), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1352]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__73_ ( .D(aes_core_keymem_n1500), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1353]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__74_ ( .D(aes_core_keymem_n1488), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1354]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__75_ ( .D(aes_core_keymem_n1476), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1355]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__76_ ( .D(aes_core_keymem_n1464), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1356]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__77_ ( .D(aes_core_keymem_n1452), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1357]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__78_ ( .D(aes_core_keymem_n1440), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1358]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__79_ ( .D(aes_core_keymem_n1428), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1359]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__80_ ( .D(aes_core_keymem_n1416), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1360]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__81_ ( .D(aes_core_keymem_n1404), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1361]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__82_ ( .D(aes_core_keymem_n1392), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1362]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__83_ ( .D(aes_core_keymem_n1380), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1363]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__84_ ( .D(aes_core_keymem_n1368), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1364]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__85_ ( .D(aes_core_keymem_n1356), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1365]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__86_ ( .D(aes_core_keymem_n1344), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1366]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__87_ ( .D(aes_core_keymem_n1332), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1367]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__88_ ( .D(aes_core_keymem_n1320), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1368]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__89_ ( .D(aes_core_keymem_n1308), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1369]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__90_ ( .D(aes_core_keymem_n1296), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1370]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__91_ ( .D(aes_core_keymem_n1284), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1371]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__92_ ( .D(aes_core_keymem_n1272), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1372]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__93_ ( .D(aes_core_keymem_n1260), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1373]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__94_ ( .D(aes_core_keymem_n1248), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1374]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__95_ ( .D(aes_core_keymem_n1236), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1375]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__96_ ( .D(aes_core_keymem_n1224), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1376]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__97_ ( .D(aes_core_keymem_n1212), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1377]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__98_ ( .D(aes_core_keymem_n1200), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1378]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__99_ ( .D(aes_core_keymem_n1188), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1379]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__100_ ( .D(aes_core_keymem_n1176), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1380]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__101_ ( .D(aes_core_keymem_n1164), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1381]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__102_ ( .D(aes_core_keymem_n1152), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1382]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__103_ ( .D(aes_core_keymem_n1140), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1383]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__104_ ( .D(aes_core_keymem_n1128), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1384]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__105_ ( .D(aes_core_keymem_n1116), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1385]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__106_ ( .D(aes_core_keymem_n1104), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1386]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__107_ ( .D(aes_core_keymem_n1092), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1387]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__108_ ( .D(aes_core_keymem_n1080), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1388]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__109_ ( .D(aes_core_keymem_n1068), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1389]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__110_ ( .D(aes_core_keymem_n1056), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1390]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__111_ ( .D(aes_core_keymem_n1044), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1391]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__112_ ( .D(aes_core_keymem_n1032), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1392]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__113_ ( .D(aes_core_keymem_n1020), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1393]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__114_ ( .D(aes_core_keymem_n1008), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1394]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__115_ ( .D(aes_core_keymem_n996), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1395]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__116_ ( .D(aes_core_keymem_n984), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1396]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__117_ ( .D(aes_core_keymem_n972), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1397]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__118_ ( .D(aes_core_keymem_n960), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1398]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__119_ ( .D(aes_core_keymem_n948), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1399]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__120_ ( .D(aes_core_keymem_n936), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1400]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__121_ ( .D(aes_core_keymem_n924), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1401]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__122_ ( .D(aes_core_keymem_n912), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1402]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__123_ ( .D(aes_core_keymem_n900), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1403]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__124_ ( .D(aes_core_keymem_n888), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1404]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__125_ ( .D(aes_core_keymem_n876), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1405]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__126_ ( .D(aes_core_keymem_n864), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1406]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_0__127_ ( .D(aes_core_keymem_n852), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1407]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__0_ ( .D(aes_core_keymem_n2374), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1024]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__8_ ( .D(aes_core_keymem_n2278), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1032]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__9_ ( .D(aes_core_keymem_n2266), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1033]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__10_ ( .D(aes_core_keymem_n2254), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1034]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__11_ ( .D(aes_core_keymem_n2242), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1035]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__12_ ( .D(aes_core_keymem_n2230), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1036]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__13_ ( .D(aes_core_keymem_n2218), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1037]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__14_ ( .D(aes_core_keymem_n2206), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1038]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__15_ ( .D(aes_core_keymem_n2194), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1039]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__16_ ( .D(aes_core_keymem_n2182), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1040]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__24_ ( .D(aes_core_keymem_n2086), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1048]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__25_ ( .D(aes_core_keymem_n2074), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1049]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__26_ ( .D(aes_core_keymem_n2062), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1050]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__27_ ( .D(aes_core_keymem_n2050), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1051]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__28_ ( .D(aes_core_keymem_n2038), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1052]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__29_ ( .D(aes_core_keymem_n2026), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1053]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__30_ ( .D(aes_core_keymem_n2014), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1054]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__31_ ( .D(aes_core_keymem_n2002), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1055]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__32_ ( .D(aes_core_keymem_n1990), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1056]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__40_ ( .D(aes_core_keymem_n1894), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1064]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__41_ ( .D(aes_core_keymem_n1882), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1065]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__42_ ( .D(aes_core_keymem_n1870), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1066]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__43_ ( .D(aes_core_keymem_n1858), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1067]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__44_ ( .D(aes_core_keymem_n1846), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1068]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__45_ ( .D(aes_core_keymem_n1834), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1069]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__46_ ( .D(aes_core_keymem_n1822), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1070]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__47_ ( .D(aes_core_keymem_n1810), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1071]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__48_ ( .D(aes_core_keymem_n1798), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1072]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__56_ ( .D(aes_core_keymem_n1702), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1080]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__57_ ( .D(aes_core_keymem_n1690), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1081]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__58_ ( .D(aes_core_keymem_n1678), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1082]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__59_ ( .D(aes_core_keymem_n1666), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1083]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__60_ ( .D(aes_core_keymem_n1654), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1084]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__61_ ( .D(aes_core_keymem_n1642), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1085]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__62_ ( .D(aes_core_keymem_n1630), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1086]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__63_ ( .D(aes_core_keymem_n1618), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1087]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__64_ ( .D(aes_core_keymem_n1606), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1088]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__72_ ( .D(aes_core_keymem_n1510), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1096]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__73_ ( .D(aes_core_keymem_n1498), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1097]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__74_ ( .D(aes_core_keymem_n1486), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1098]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__75_ ( .D(aes_core_keymem_n1474), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1099]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__76_ ( .D(aes_core_keymem_n1462), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1100]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__77_ ( .D(aes_core_keymem_n1450), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1101]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__78_ ( .D(aes_core_keymem_n1438), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1102]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__79_ ( .D(aes_core_keymem_n1426), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1103]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__80_ ( .D(aes_core_keymem_n1414), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1104]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__88_ ( .D(aes_core_keymem_n1318), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1112]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__89_ ( .D(aes_core_keymem_n1306), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1113]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__90_ ( .D(aes_core_keymem_n1294), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1114]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__91_ ( .D(aes_core_keymem_n1282), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1115]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__92_ ( .D(aes_core_keymem_n1270), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1116]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__93_ ( .D(aes_core_keymem_n1258), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1117]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__94_ ( .D(aes_core_keymem_n1246), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1118]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__95_ ( .D(aes_core_keymem_n1234), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1119]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__96_ ( .D(aes_core_keymem_n1222), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1120]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__104_ ( .D(aes_core_keymem_n1126), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1128]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__105_ ( .D(aes_core_keymem_n1114), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1129]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__106_ ( .D(aes_core_keymem_n1102), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1130]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__107_ ( .D(aes_core_keymem_n1090), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1131]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__108_ ( .D(aes_core_keymem_n1078), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1132]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__109_ ( .D(aes_core_keymem_n1066), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1133]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__110_ ( .D(aes_core_keymem_n1054), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1134]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__111_ ( .D(aes_core_keymem_n1042), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1135]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__112_ ( .D(aes_core_keymem_n1030), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1136]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__120_ ( .D(aes_core_keymem_n934), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1144]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__121_ ( .D(aes_core_keymem_n922), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1145]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__122_ ( .D(aes_core_keymem_n910), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1146]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__123_ ( .D(aes_core_keymem_n898), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1147]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__124_ ( .D(aes_core_keymem_n886), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1148]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__125_ ( .D(aes_core_keymem_n874), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1149]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__126_ ( .D(aes_core_keymem_n862), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1150]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_2__127_ ( .D(aes_core_keymem_n850), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1151]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__0_ ( .D(aes_core_keymem_n2373), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[896]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__8_ ( .D(aes_core_keymem_n2277), .CK(
        clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[904]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__10_ ( .D(aes_core_keymem_n2253), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[906]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__13_ ( .D(aes_core_keymem_n2217), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[909]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__14_ ( .D(aes_core_keymem_n2205), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[910]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__15_ ( .D(aes_core_keymem_n2193), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[911]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__16_ ( .D(aes_core_keymem_n2181), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[912]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__24_ ( .D(aes_core_keymem_n2085), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[920]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__26_ ( .D(aes_core_keymem_n2061), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[922]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__29_ ( .D(aes_core_keymem_n2025), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[925]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__30_ ( .D(aes_core_keymem_n2013), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[926]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__31_ ( .D(aes_core_keymem_n2001), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[927]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__32_ ( .D(aes_core_keymem_n1989), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[928]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__40_ ( .D(aes_core_keymem_n1893), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[936]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__42_ ( .D(aes_core_keymem_n1869), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[938]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__45_ ( .D(aes_core_keymem_n1833), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[941]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__46_ ( .D(aes_core_keymem_n1821), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[942]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__47_ ( .D(aes_core_keymem_n1809), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[943]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__48_ ( .D(aes_core_keymem_n1797), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[944]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__56_ ( .D(aes_core_keymem_n1701), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[952]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__58_ ( .D(aes_core_keymem_n1677), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[954]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__61_ ( .D(aes_core_keymem_n1641), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[957]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__62_ ( .D(aes_core_keymem_n1629), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[958]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__63_ ( .D(aes_core_keymem_n1617), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[959]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__64_ ( .D(aes_core_keymem_n1605), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[960]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__72_ ( .D(aes_core_keymem_n1509), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[968]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__74_ ( .D(aes_core_keymem_n1485), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[970]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__77_ ( .D(aes_core_keymem_n1449), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[973]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__78_ ( .D(aes_core_keymem_n1437), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[974]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__79_ ( .D(aes_core_keymem_n1425), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[975]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__80_ ( .D(aes_core_keymem_n1413), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[976]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__88_ ( .D(aes_core_keymem_n1317), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[984]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__90_ ( .D(aes_core_keymem_n1293), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[986]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__93_ ( .D(aes_core_keymem_n1257), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[989]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__94_ ( .D(aes_core_keymem_n1245), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[990]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__95_ ( .D(aes_core_keymem_n1233), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[991]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__96_ ( .D(aes_core_keymem_n1221), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[992]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__104_ ( .D(aes_core_keymem_n1125), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1000]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__106_ ( .D(aes_core_keymem_n1101), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1002]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__109_ ( .D(aes_core_keymem_n1065), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1005]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__110_ ( .D(aes_core_keymem_n1053), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1006]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__111_ ( .D(aes_core_keymem_n1041), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1007]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__112_ ( .D(aes_core_keymem_n1029), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1008]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__120_ ( .D(aes_core_keymem_n933), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1016]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__122_ ( .D(aes_core_keymem_n909), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1018]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__125_ ( .D(aes_core_keymem_n873), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1021]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__126_ ( .D(aes_core_keymem_n861), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1022]) );
  DFFRHQX1 aes_core_keymem_key_mem_reg_3__127_ ( .D(aes_core_keymem_n849), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem[1023]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_32_ ( .D(aes_core_keymem_n1993), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[32]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_33_ ( .D(aes_core_keymem_n1981), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[33]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_34_ ( .D(aes_core_keymem_n1969), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[34]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_35_ ( .D(aes_core_keymem_n1957), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[35]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_36_ ( .D(aes_core_keymem_n1945), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[36]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_37_ ( .D(aes_core_keymem_n1933), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[37]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_38_ ( .D(aes_core_keymem_n1921), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[38]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_39_ ( .D(aes_core_keymem_n1909), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[39]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_40_ ( .D(aes_core_keymem_n1897), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[40]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_41_ ( .D(aes_core_keymem_n1885), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[41]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_42_ ( .D(aes_core_keymem_n1873), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[42]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_43_ ( .D(aes_core_keymem_n1861), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[43]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_44_ ( .D(aes_core_keymem_n1849), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[44]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_45_ ( .D(aes_core_keymem_n1837), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[45]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_46_ ( .D(aes_core_keymem_n1825), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[46]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_47_ ( .D(aes_core_keymem_n1813), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[47]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_48_ ( .D(aes_core_keymem_n1801), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[48]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_49_ ( .D(aes_core_keymem_n1789), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[49]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_50_ ( .D(aes_core_keymem_n1777), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[50]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_51_ ( .D(aes_core_keymem_n1765), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[51]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_52_ ( .D(aes_core_keymem_n1753), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[52]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_53_ ( .D(aes_core_keymem_n1741), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[53]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_54_ ( .D(aes_core_keymem_n1729), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[54]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_55_ ( .D(aes_core_keymem_n1717), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[55]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_56_ ( .D(aes_core_keymem_n1705), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[56]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_57_ ( .D(aes_core_keymem_n1693), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[57]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_58_ ( .D(aes_core_keymem_n1681), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[58]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_59_ ( .D(aes_core_keymem_n1669), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[59]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_60_ ( .D(aes_core_keymem_n1657), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[60]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_61_ ( .D(aes_core_keymem_n1645), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[61]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_62_ ( .D(aes_core_keymem_n1633), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[62]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_63_ ( .D(aes_core_keymem_n1621), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[63]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_64_ ( .D(aes_core_keymem_n1609), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[64]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_65_ ( .D(aes_core_keymem_n1597), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[65]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_66_ ( .D(aes_core_keymem_n1585), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[66]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_67_ ( .D(aes_core_keymem_n1573), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[67]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_68_ ( .D(aes_core_keymem_n1561), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[68]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_69_ ( .D(aes_core_keymem_n1549), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[69]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_70_ ( .D(aes_core_keymem_n1537), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[70]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_71_ ( .D(aes_core_keymem_n1525), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[71]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_72_ ( .D(aes_core_keymem_n1513), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[72]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_73_ ( .D(aes_core_keymem_n1501), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[73]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_74_ ( .D(aes_core_keymem_n1489), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[74]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_75_ ( .D(aes_core_keymem_n1477), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[75]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_76_ ( .D(aes_core_keymem_n1465), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[76]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_77_ ( .D(aes_core_keymem_n1453), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[77]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_78_ ( .D(aes_core_keymem_n1441), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[78]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_79_ ( .D(aes_core_keymem_n1429), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[79]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_80_ ( .D(aes_core_keymem_n1417), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[80]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_81_ ( .D(aes_core_keymem_n1405), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[81]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_82_ ( .D(aes_core_keymem_n1393), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[82]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_83_ ( .D(aes_core_keymem_n1381), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[83]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_84_ ( .D(aes_core_keymem_n1369), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[84]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_85_ ( .D(aes_core_keymem_n1357), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[85]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_86_ ( .D(aes_core_keymem_n1345), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[86]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_87_ ( .D(aes_core_keymem_n1333), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[87]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_88_ ( .D(aes_core_keymem_n1321), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[88]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_89_ ( .D(aes_core_keymem_n1309), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[89]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_90_ ( .D(aes_core_keymem_n1297), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[90]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_91_ ( .D(aes_core_keymem_n1285), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[91]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_92_ ( .D(aes_core_keymem_n1273), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[92]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_93_ ( .D(aes_core_keymem_n1261), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[93]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_94_ ( .D(aes_core_keymem_n1249), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[94]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_95_ ( .D(aes_core_keymem_n1237), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[95]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_96_ ( .D(aes_core_keymem_n1225), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[96]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_97_ ( .D(aes_core_keymem_n1213), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[97]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_98_ ( .D(aes_core_keymem_n1201), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[98]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_99_ ( .D(aes_core_keymem_n1189), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[99]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_100_ ( .D(aes_core_keymem_n1177), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[100]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_101_ ( .D(aes_core_keymem_n1165), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[101]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_102_ ( .D(aes_core_keymem_n1153), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[102]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_103_ ( .D(aes_core_keymem_n1141), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[103]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_104_ ( .D(aes_core_keymem_n1129), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[104]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_105_ ( .D(aes_core_keymem_n1117), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[105]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_106_ ( .D(aes_core_keymem_n1105), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[106]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_107_ ( .D(aes_core_keymem_n1093), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[107]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_108_ ( .D(aes_core_keymem_n1081), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[108]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_109_ ( .D(aes_core_keymem_n1069), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[109]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_110_ ( .D(aes_core_keymem_n1057), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[110]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_111_ ( .D(aes_core_keymem_n1045), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[111]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_112_ ( .D(aes_core_keymem_n1033), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[112]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_113_ ( .D(aes_core_keymem_n1021), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[113]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_114_ ( .D(aes_core_keymem_n1009), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[114]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_115_ ( .D(aes_core_keymem_n997), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[115]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_116_ ( .D(aes_core_keymem_n985), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[116]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_117_ ( .D(aes_core_keymem_n973), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[117]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_118_ ( .D(aes_core_keymem_n961), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[118]) );
  DFFHQX1 aes_core_keymem_prev_key1_reg_reg_119_ ( .D(aes_core_keymem_n949), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_prev_key1_reg[119]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__0_ ( .D(aes_core_keymem_n2371), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[256]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__1_ ( .D(aes_core_keymem_n2359), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[257]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__2_ ( .D(aes_core_keymem_n2347), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[258]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__3_ ( .D(aes_core_keymem_n2335), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[259]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__4_ ( .D(aes_core_keymem_n2323), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[260]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__5_ ( .D(aes_core_keymem_n2311), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[261]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__6_ ( .D(aes_core_keymem_n2299), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[262]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__7_ ( .D(aes_core_keymem_n2287), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[263]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__8_ ( .D(aes_core_keymem_n2275), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[264]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__9_ ( .D(aes_core_keymem_n2263), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[265]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__10_ ( .D(aes_core_keymem_n2251), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[266]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__11_ ( .D(aes_core_keymem_n2239), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[267]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__12_ ( .D(aes_core_keymem_n2227), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[268]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__13_ ( .D(aes_core_keymem_n2215), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[269]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__14_ ( .D(aes_core_keymem_n2203), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[270]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__15_ ( .D(aes_core_keymem_n2191), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[271]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__16_ ( .D(aes_core_keymem_n2179), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[272]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__17_ ( .D(aes_core_keymem_n2167), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[273]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__18_ ( .D(aes_core_keymem_n2155), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[274]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__19_ ( .D(aes_core_keymem_n2143), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[275]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__20_ ( .D(aes_core_keymem_n2131), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[276]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__21_ ( .D(aes_core_keymem_n2119), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[277]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__22_ ( .D(aes_core_keymem_n2107), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[278]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__23_ ( .D(aes_core_keymem_n2095), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[279]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__24_ ( .D(aes_core_keymem_n2083), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[280]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__25_ ( .D(aes_core_keymem_n2071), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[281]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__26_ ( .D(aes_core_keymem_n2059), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[282]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__27_ ( .D(aes_core_keymem_n2047), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[283]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__28_ ( .D(aes_core_keymem_n2035), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[284]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__29_ ( .D(aes_core_keymem_n2023), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[285]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__30_ ( .D(aes_core_keymem_n2011), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[286]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__31_ ( .D(aes_core_keymem_n1999), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[287]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__32_ ( .D(aes_core_keymem_n1987), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[288]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__33_ ( .D(aes_core_keymem_n1975), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[289]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__34_ ( .D(aes_core_keymem_n1963), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[290]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__35_ ( .D(aes_core_keymem_n1951), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[291]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__36_ ( .D(aes_core_keymem_n1939), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[292]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__37_ ( .D(aes_core_keymem_n1927), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[293]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__38_ ( .D(aes_core_keymem_n1915), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[294]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__39_ ( .D(aes_core_keymem_n1903), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[295]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__40_ ( .D(aes_core_keymem_n1891), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[296]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__41_ ( .D(aes_core_keymem_n1879), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[297]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__42_ ( .D(aes_core_keymem_n1867), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[298]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__43_ ( .D(aes_core_keymem_n1855), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[299]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__44_ ( .D(aes_core_keymem_n1843), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[300]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__45_ ( .D(aes_core_keymem_n1831), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[301]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__46_ ( .D(aes_core_keymem_n1819), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[302]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__47_ ( .D(aes_core_keymem_n1807), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[303]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__48_ ( .D(aes_core_keymem_n1795), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[304]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__49_ ( .D(aes_core_keymem_n1783), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[305]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__50_ ( .D(aes_core_keymem_n1771), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[306]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__51_ ( .D(aes_core_keymem_n1759), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[307]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__52_ ( .D(aes_core_keymem_n1747), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[308]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__53_ ( .D(aes_core_keymem_n1735), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[309]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__54_ ( .D(aes_core_keymem_n1723), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[310]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__55_ ( .D(aes_core_keymem_n1711), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[311]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__56_ ( .D(aes_core_keymem_n1699), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[312]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__57_ ( .D(aes_core_keymem_n1687), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[313]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__58_ ( .D(aes_core_keymem_n1675), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[314]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__59_ ( .D(aes_core_keymem_n1663), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[315]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__60_ ( .D(aes_core_keymem_n1651), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[316]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__61_ ( .D(aes_core_keymem_n1639), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[317]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__62_ ( .D(aes_core_keymem_n1627), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[318]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__63_ ( .D(aes_core_keymem_n1615), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[319]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__64_ ( .D(aes_core_keymem_n1603), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[320]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__65_ ( .D(aes_core_keymem_n1591), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[321]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__66_ ( .D(aes_core_keymem_n1579), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[322]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__67_ ( .D(aes_core_keymem_n1567), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[323]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__68_ ( .D(aes_core_keymem_n1555), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[324]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__69_ ( .D(aes_core_keymem_n1543), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[325]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__70_ ( .D(aes_core_keymem_n1531), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[326]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__71_ ( .D(aes_core_keymem_n1519), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[327]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__72_ ( .D(aes_core_keymem_n1507), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[328]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__73_ ( .D(aes_core_keymem_n1495), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[329]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__74_ ( .D(aes_core_keymem_n1483), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[330]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__75_ ( .D(aes_core_keymem_n1471), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[331]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__76_ ( .D(aes_core_keymem_n1459), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[332]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__77_ ( .D(aes_core_keymem_n1447), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[333]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__78_ ( .D(aes_core_keymem_n1435), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[334]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__79_ ( .D(aes_core_keymem_n1423), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[335]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__80_ ( .D(aes_core_keymem_n1411), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[336]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__81_ ( .D(aes_core_keymem_n1399), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[337]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__82_ ( .D(aes_core_keymem_n1387), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[338]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__83_ ( .D(aes_core_keymem_n1375), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[339]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__84_ ( .D(aes_core_keymem_n1363), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[340]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__85_ ( .D(aes_core_keymem_n1351), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[341]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__86_ ( .D(aes_core_keymem_n1339), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[342]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__87_ ( .D(aes_core_keymem_n1327), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[343]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__88_ ( .D(aes_core_keymem_n1315), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[344]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__89_ ( .D(aes_core_keymem_n1303), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[345]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__90_ ( .D(aes_core_keymem_n1291), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[346]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__91_ ( .D(aes_core_keymem_n1279), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[347]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__92_ ( .D(aes_core_keymem_n1267), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[348]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__93_ ( .D(aes_core_keymem_n1255), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[349]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__94_ ( .D(aes_core_keymem_n1243), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[350]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__95_ ( .D(aes_core_keymem_n1231), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[351]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__96_ ( .D(aes_core_keymem_n1219), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[352]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__97_ ( .D(aes_core_keymem_n1207), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[353]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__98_ ( .D(aes_core_keymem_n1195), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[354]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__99_ ( .D(aes_core_keymem_n1183), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[355]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__100_ ( .D(aes_core_keymem_n1171), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[356]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__101_ ( .D(aes_core_keymem_n1159), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[357]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__102_ ( .D(aes_core_keymem_n1147), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[358]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__103_ ( .D(aes_core_keymem_n1135), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[359]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__104_ ( .D(aes_core_keymem_n1123), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[360]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__105_ ( .D(aes_core_keymem_n1111), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[361]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__106_ ( .D(aes_core_keymem_n1099), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[362]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__107_ ( .D(aes_core_keymem_n1087), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[363]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__108_ ( .D(aes_core_keymem_n1075), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[364]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__109_ ( .D(aes_core_keymem_n1063), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[365]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__110_ ( .D(aes_core_keymem_n1051), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[366]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__111_ ( .D(aes_core_keymem_n1039), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[367]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__112_ ( .D(aes_core_keymem_n1027), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[368]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__113_ ( .D(aes_core_keymem_n1015), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[369]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__114_ ( .D(aes_core_keymem_n1003), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[370]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__115_ ( .D(aes_core_keymem_n991), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[371]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__116_ ( .D(aes_core_keymem_n979), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[372]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__117_ ( .D(aes_core_keymem_n967), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[373]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__118_ ( .D(aes_core_keymem_n955), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[374]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__119_ ( .D(aes_core_keymem_n943), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[375]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__120_ ( .D(aes_core_keymem_n931), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[376]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__121_ ( .D(aes_core_keymem_n919), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[377]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__122_ ( .D(aes_core_keymem_n907), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[378]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__123_ ( .D(aes_core_keymem_n895), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[379]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__124_ ( .D(aes_core_keymem_n883), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[380]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__125_ ( .D(aes_core_keymem_n871), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[381]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__126_ ( .D(aes_core_keymem_n859), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[382]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_5__127_ ( .D(aes_core_keymem_n847), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[383]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__0_ ( .D(aes_core_keymem_n2368), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[768]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__1_ ( .D(aes_core_keymem_n2356), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[769]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__2_ ( .D(aes_core_keymem_n2344), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[770]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__3_ ( .D(aes_core_keymem_n2332), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[771]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__4_ ( .D(aes_core_keymem_n2320), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[772]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__5_ ( .D(aes_core_keymem_n2308), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[773]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__6_ ( .D(aes_core_keymem_n2296), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[774]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__7_ ( .D(aes_core_keymem_n2284), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[775]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__8_ ( .D(aes_core_keymem_n2272), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[776]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__9_ ( .D(aes_core_keymem_n2260), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[777]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__10_ ( .D(aes_core_keymem_n2248), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[778]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__11_ ( .D(aes_core_keymem_n2236), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[779]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__12_ ( .D(aes_core_keymem_n2224), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[780]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__13_ ( .D(aes_core_keymem_n2212), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[781]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__14_ ( .D(aes_core_keymem_n2200), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[782]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__15_ ( .D(aes_core_keymem_n2188), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[783]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__16_ ( .D(aes_core_keymem_n2176), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[784]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__17_ ( .D(aes_core_keymem_n2164), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[785]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__18_ ( .D(aes_core_keymem_n2152), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[786]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__19_ ( .D(aes_core_keymem_n2140), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[787]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__20_ ( .D(aes_core_keymem_n2128), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[788]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__21_ ( .D(aes_core_keymem_n2116), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[789]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__22_ ( .D(aes_core_keymem_n2104), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[790]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__23_ ( .D(aes_core_keymem_n2092), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[791]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__24_ ( .D(aes_core_keymem_n2080), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[792]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__25_ ( .D(aes_core_keymem_n2068), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[793]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__26_ ( .D(aes_core_keymem_n2056), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[794]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__27_ ( .D(aes_core_keymem_n2044), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[795]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__28_ ( .D(aes_core_keymem_n2032), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[796]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__29_ ( .D(aes_core_keymem_n2020), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[797]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__30_ ( .D(aes_core_keymem_n2008), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[798]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__31_ ( .D(aes_core_keymem_n1996), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[799]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__32_ ( .D(aes_core_keymem_n1984), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[800]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__33_ ( .D(aes_core_keymem_n1972), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[801]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__34_ ( .D(aes_core_keymem_n1960), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[802]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__35_ ( .D(aes_core_keymem_n1948), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[803]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__36_ ( .D(aes_core_keymem_n1936), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[804]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__37_ ( .D(aes_core_keymem_n1924), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[805]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__38_ ( .D(aes_core_keymem_n1912), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[806]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__39_ ( .D(aes_core_keymem_n1900), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[807]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__40_ ( .D(aes_core_keymem_n1888), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[808]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__41_ ( .D(aes_core_keymem_n1876), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[809]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__42_ ( .D(aes_core_keymem_n1864), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[810]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__43_ ( .D(aes_core_keymem_n1852), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[811]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__44_ ( .D(aes_core_keymem_n1840), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[812]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__45_ ( .D(aes_core_keymem_n1828), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[813]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__46_ ( .D(aes_core_keymem_n1816), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[814]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__47_ ( .D(aes_core_keymem_n1804), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[815]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__48_ ( .D(aes_core_keymem_n1792), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[816]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__49_ ( .D(aes_core_keymem_n1780), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[817]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__50_ ( .D(aes_core_keymem_n1768), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[818]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__51_ ( .D(aes_core_keymem_n1756), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[819]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__52_ ( .D(aes_core_keymem_n1744), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[820]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__53_ ( .D(aes_core_keymem_n1732), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[821]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__54_ ( .D(aes_core_keymem_n1720), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[822]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__55_ ( .D(aes_core_keymem_n1708), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[823]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__56_ ( .D(aes_core_keymem_n1696), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[824]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__57_ ( .D(aes_core_keymem_n1684), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[825]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__58_ ( .D(aes_core_keymem_n1672), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[826]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__59_ ( .D(aes_core_keymem_n1660), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[827]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__60_ ( .D(aes_core_keymem_n1648), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[828]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__61_ ( .D(aes_core_keymem_n1636), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[829]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__62_ ( .D(aes_core_keymem_n1624), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[830]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__63_ ( .D(aes_core_keymem_n1612), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[831]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__64_ ( .D(aes_core_keymem_n1600), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[832]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__65_ ( .D(aes_core_keymem_n1588), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[833]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__66_ ( .D(aes_core_keymem_n1576), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[834]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__67_ ( .D(aes_core_keymem_n1564), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[835]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__68_ ( .D(aes_core_keymem_n1552), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[836]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__69_ ( .D(aes_core_keymem_n1540), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[837]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__70_ ( .D(aes_core_keymem_n1528), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[838]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__71_ ( .D(aes_core_keymem_n1516), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[839]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__72_ ( .D(aes_core_keymem_n1504), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[840]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__73_ ( .D(aes_core_keymem_n1492), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[841]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__74_ ( .D(aes_core_keymem_n1480), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[842]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__75_ ( .D(aes_core_keymem_n1468), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[843]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__76_ ( .D(aes_core_keymem_n1456), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[844]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__77_ ( .D(aes_core_keymem_n1444), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[845]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__78_ ( .D(aes_core_keymem_n1432), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[846]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__79_ ( .D(aes_core_keymem_n1420), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[847]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__80_ ( .D(aes_core_keymem_n1408), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[848]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__81_ ( .D(aes_core_keymem_n1396), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[849]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__82_ ( .D(aes_core_keymem_n1384), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[850]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__83_ ( .D(aes_core_keymem_n1372), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[851]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__84_ ( .D(aes_core_keymem_n1360), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[852]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__85_ ( .D(aes_core_keymem_n1348), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[853]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__86_ ( .D(aes_core_keymem_n1336), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[854]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__87_ ( .D(aes_core_keymem_n1324), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[855]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__88_ ( .D(aes_core_keymem_n1312), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[856]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__89_ ( .D(aes_core_keymem_n1300), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[857]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__90_ ( .D(aes_core_keymem_n1288), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[858]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__91_ ( .D(aes_core_keymem_n1276), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[859]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__92_ ( .D(aes_core_keymem_n1264), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[860]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__93_ ( .D(aes_core_keymem_n1252), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[861]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__94_ ( .D(aes_core_keymem_n1240), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[862]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__95_ ( .D(aes_core_keymem_n1228), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[863]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__96_ ( .D(aes_core_keymem_n1216), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[864]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__97_ ( .D(aes_core_keymem_n1204), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[865]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__98_ ( .D(aes_core_keymem_n1192), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[866]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__99_ ( .D(aes_core_keymem_n1180), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[867]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__100_ ( .D(aes_core_keymem_n1168), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[868]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__101_ ( .D(aes_core_keymem_n1156), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[869]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__102_ ( .D(aes_core_keymem_n1144), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[870]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__103_ ( .D(aes_core_keymem_n1132), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[871]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__104_ ( .D(aes_core_keymem_n1120), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[872]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__105_ ( .D(aes_core_keymem_n1108), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[873]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__106_ ( .D(aes_core_keymem_n1096), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[874]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__107_ ( .D(aes_core_keymem_n1084), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[875]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__108_ ( .D(aes_core_keymem_n1072), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[876]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__109_ ( .D(aes_core_keymem_n1060), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[877]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__110_ ( .D(aes_core_keymem_n1048), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[878]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__111_ ( .D(aes_core_keymem_n1036), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[879]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__112_ ( .D(aes_core_keymem_n1024), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[880]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__113_ ( .D(aes_core_keymem_n1012), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[881]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__114_ ( .D(aes_core_keymem_n1000), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[882]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__115_ ( .D(aes_core_keymem_n988), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[883]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__116_ ( .D(aes_core_keymem_n976), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[884]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__117_ ( .D(aes_core_keymem_n964), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[885]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__118_ ( .D(aes_core_keymem_n952), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[886]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__119_ ( .D(aes_core_keymem_n940), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[887]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__120_ ( .D(aes_core_keymem_n928), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[888]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__121_ ( .D(aes_core_keymem_n916), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[889]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__122_ ( .D(aes_core_keymem_n904), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[890]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__123_ ( .D(aes_core_keymem_n892), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[891]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__124_ ( .D(aes_core_keymem_n880), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[892]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__125_ ( .D(aes_core_keymem_n868), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[893]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__126_ ( .D(aes_core_keymem_n856), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[894]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_8__127_ ( .D(aes_core_keymem_n844), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[895]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__0_ ( .D(aes_core_keymem_n2372), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[384]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__8_ ( .D(aes_core_keymem_n2276), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[392]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__10_ ( .D(aes_core_keymem_n2252), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[394]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__13_ ( .D(aes_core_keymem_n2216), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[397]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__14_ ( .D(aes_core_keymem_n2204), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[398]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__15_ ( .D(aes_core_keymem_n2192), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[399]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__16_ ( .D(aes_core_keymem_n2180), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[400]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__24_ ( .D(aes_core_keymem_n2084), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[408]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__25_ ( .D(aes_core_keymem_n2072), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[409]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__26_ ( .D(aes_core_keymem_n2060), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[410]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__27_ ( .D(aes_core_keymem_n2048), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[411]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__28_ ( .D(aes_core_keymem_n2036), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[412]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__29_ ( .D(aes_core_keymem_n2024), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[413]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__30_ ( .D(aes_core_keymem_n2012), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[414]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__31_ ( .D(aes_core_keymem_n2000), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[415]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__32_ ( .D(aes_core_keymem_n1988), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[416]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__40_ ( .D(aes_core_keymem_n1892), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[424]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__42_ ( .D(aes_core_keymem_n1868), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[426]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__45_ ( .D(aes_core_keymem_n1832), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[429]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__46_ ( .D(aes_core_keymem_n1820), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[430]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__47_ ( .D(aes_core_keymem_n1808), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[431]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__48_ ( .D(aes_core_keymem_n1796), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[432]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__56_ ( .D(aes_core_keymem_n1700), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[440]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__57_ ( .D(aes_core_keymem_n1688), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[441]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__58_ ( .D(aes_core_keymem_n1676), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[442]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__59_ ( .D(aes_core_keymem_n1664), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[443]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__60_ ( .D(aes_core_keymem_n1652), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[444]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__61_ ( .D(aes_core_keymem_n1640), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[445]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__62_ ( .D(aes_core_keymem_n1628), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[446]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__63_ ( .D(aes_core_keymem_n1616), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[447]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__64_ ( .D(aes_core_keymem_n1604), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[448]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__72_ ( .D(aes_core_keymem_n1508), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[456]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__74_ ( .D(aes_core_keymem_n1484), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[458]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__77_ ( .D(aes_core_keymem_n1448), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[461]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__78_ ( .D(aes_core_keymem_n1436), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[462]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__79_ ( .D(aes_core_keymem_n1424), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[463]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__80_ ( .D(aes_core_keymem_n1412), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[464]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__88_ ( .D(aes_core_keymem_n1316), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[472]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__89_ ( .D(aes_core_keymem_n1304), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[473]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__90_ ( .D(aes_core_keymem_n1292), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[474]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__91_ ( .D(aes_core_keymem_n1280), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[475]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__92_ ( .D(aes_core_keymem_n1268), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[476]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__93_ ( .D(aes_core_keymem_n1256), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[477]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__94_ ( .D(aes_core_keymem_n1244), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[478]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__95_ ( .D(aes_core_keymem_n1232), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[479]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__96_ ( .D(aes_core_keymem_n1220), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[480]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__104_ ( .D(aes_core_keymem_n1124), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[488]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__106_ ( .D(aes_core_keymem_n1100), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[490]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__109_ ( .D(aes_core_keymem_n1064), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[493]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__110_ ( .D(aes_core_keymem_n1052), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[494]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__111_ ( .D(aes_core_keymem_n1040), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[495]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__112_ ( .D(aes_core_keymem_n1028), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[496]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__120_ ( .D(aes_core_keymem_n932), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[504]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__121_ ( .D(aes_core_keymem_n920), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[505]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__122_ ( .D(aes_core_keymem_n908), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[506]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__123_ ( .D(aes_core_keymem_n896), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[507]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__124_ ( .D(aes_core_keymem_n884), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[508]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__125_ ( .D(aes_core_keymem_n872), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[509]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__126_ ( .D(aes_core_keymem_n860), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[510]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_4__127_ ( .D(aes_core_keymem_n848), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[511]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__0_ ( .D(aes_core_keymem_n2369), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[0]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__8_ ( .D(aes_core_keymem_n2273), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[8]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__10_ ( .D(aes_core_keymem_n2249), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[10]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__13_ ( .D(aes_core_keymem_n2213), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[13]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__14_ ( .D(aes_core_keymem_n2201), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[14]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__15_ ( .D(aes_core_keymem_n2189), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[15]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__16_ ( .D(aes_core_keymem_n2177), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[16]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__24_ ( .D(aes_core_keymem_n2081), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[24]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__25_ ( .D(aes_core_keymem_n2069), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[25]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__26_ ( .D(aes_core_keymem_n2057), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[26]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__27_ ( .D(aes_core_keymem_n2045), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[27]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__28_ ( .D(aes_core_keymem_n2033), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[28]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__29_ ( .D(aes_core_keymem_n2021), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[29]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__30_ ( .D(aes_core_keymem_n2009), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[30]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__31_ ( .D(aes_core_keymem_n1997), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[31]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__32_ ( .D(aes_core_keymem_n1985), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[32]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__40_ ( .D(aes_core_keymem_n1889), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[40]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__42_ ( .D(aes_core_keymem_n1865), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[42]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__45_ ( .D(aes_core_keymem_n1829), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[45]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__46_ ( .D(aes_core_keymem_n1817), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[46]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__47_ ( .D(aes_core_keymem_n1805), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[47]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__48_ ( .D(aes_core_keymem_n1793), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[48]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__56_ ( .D(aes_core_keymem_n1697), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[56]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__57_ ( .D(aes_core_keymem_n1685), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[57]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__58_ ( .D(aes_core_keymem_n1673), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[58]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__59_ ( .D(aes_core_keymem_n1661), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[59]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__60_ ( .D(aes_core_keymem_n1649), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[60]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__61_ ( .D(aes_core_keymem_n1637), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[61]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__62_ ( .D(aes_core_keymem_n1625), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[62]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__63_ ( .D(aes_core_keymem_n1613), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[63]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__64_ ( .D(aes_core_keymem_n1601), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[64]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__72_ ( .D(aes_core_keymem_n1505), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[72]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__74_ ( .D(aes_core_keymem_n1481), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[74]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__77_ ( .D(aes_core_keymem_n1445), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[77]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__78_ ( .D(aes_core_keymem_n1433), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[78]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__79_ ( .D(aes_core_keymem_n1421), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[79]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__80_ ( .D(aes_core_keymem_n1409), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[80]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__88_ ( .D(aes_core_keymem_n1313), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[88]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__89_ ( .D(aes_core_keymem_n1301), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[89]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__90_ ( .D(aes_core_keymem_n1289), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[90]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__91_ ( .D(aes_core_keymem_n1277), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[91]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__92_ ( .D(aes_core_keymem_n1265), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[92]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__93_ ( .D(aes_core_keymem_n1253), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[93]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__94_ ( .D(aes_core_keymem_n1241), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[94]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__95_ ( .D(aes_core_keymem_n1229), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[95]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__96_ ( .D(aes_core_keymem_n1217), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[96]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__104_ ( .D(aes_core_keymem_n1121), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[104]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__106_ ( .D(aes_core_keymem_n1097), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[106]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__109_ ( .D(aes_core_keymem_n1061), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[109]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__110_ ( .D(aes_core_keymem_n1049), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[110]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__111_ ( .D(aes_core_keymem_n1037), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[111]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__112_ ( .D(aes_core_keymem_n1025), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[112]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__120_ ( .D(aes_core_keymem_n929), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[120]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__121_ ( .D(aes_core_keymem_n917), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[121]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__122_ ( .D(aes_core_keymem_n905), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[122]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__123_ ( .D(aes_core_keymem_n893), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[123]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__124_ ( .D(aes_core_keymem_n881), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[124]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__125_ ( .D(aes_core_keymem_n869), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[125]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__126_ ( .D(aes_core_keymem_n857), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[126]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_7__127_ ( .D(aes_core_keymem_n845), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[127]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__0_ ( .D(aes_core_keymem_n2370), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[128]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__8_ ( .D(aes_core_keymem_n2274), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[136]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__10_ ( .D(aes_core_keymem_n2250), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[138]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__13_ ( .D(aes_core_keymem_n2214), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[141]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__14_ ( .D(aes_core_keymem_n2202), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[142]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__15_ ( .D(aes_core_keymem_n2190), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[143]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__16_ ( .D(aes_core_keymem_n2178), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[144]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__24_ ( .D(aes_core_keymem_n2082), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[152]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__26_ ( .D(aes_core_keymem_n2058), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[154]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__29_ ( .D(aes_core_keymem_n2022), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[157]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__30_ ( .D(aes_core_keymem_n2010), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[158]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__31_ ( .D(aes_core_keymem_n1998), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[159]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__32_ ( .D(aes_core_keymem_n1986), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[160]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__40_ ( .D(aes_core_keymem_n1890), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[168]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__42_ ( .D(aes_core_keymem_n1866), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[170]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__45_ ( .D(aes_core_keymem_n1830), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[173]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__46_ ( .D(aes_core_keymem_n1818), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[174]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__47_ ( .D(aes_core_keymem_n1806), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[175]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__48_ ( .D(aes_core_keymem_n1794), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[176]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__56_ ( .D(aes_core_keymem_n1698), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[184]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__58_ ( .D(aes_core_keymem_n1674), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[186]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__61_ ( .D(aes_core_keymem_n1638), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[189]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__62_ ( .D(aes_core_keymem_n1626), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[190]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__63_ ( .D(aes_core_keymem_n1614), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[191]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__64_ ( .D(aes_core_keymem_n1602), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[192]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__72_ ( .D(aes_core_keymem_n1506), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[200]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__74_ ( .D(aes_core_keymem_n1482), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[202]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__77_ ( .D(aes_core_keymem_n1446), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[205]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__78_ ( .D(aes_core_keymem_n1434), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[206]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__79_ ( .D(aes_core_keymem_n1422), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[207]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__80_ ( .D(aes_core_keymem_n1410), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[208]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__88_ ( .D(aes_core_keymem_n1314), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[216]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__90_ ( .D(aes_core_keymem_n1290), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[218]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__93_ ( .D(aes_core_keymem_n1254), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[221]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__94_ ( .D(aes_core_keymem_n1242), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[222]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__95_ ( .D(aes_core_keymem_n1230), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[223]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__96_ ( .D(aes_core_keymem_n1218), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[224]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__104_ ( .D(aes_core_keymem_n1122), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[232]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__106_ ( .D(aes_core_keymem_n1098), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[234]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__109_ ( .D(aes_core_keymem_n1062), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[237]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__110_ ( .D(aes_core_keymem_n1050), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[238]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__111_ ( .D(aes_core_keymem_n1038), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[239]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__112_ ( .D(aes_core_keymem_n1026), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[240]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__120_ ( .D(aes_core_keymem_n930), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[248]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__122_ ( .D(aes_core_keymem_n906), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[250]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__125_ ( .D(aes_core_keymem_n870), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[253]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__126_ ( .D(aes_core_keymem_n858), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[254]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_6__127_ ( .D(aes_core_keymem_n846), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[255]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__0_ ( .D(aes_core_keymem_n2367), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[640]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__8_ ( .D(aes_core_keymem_n2271), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[648]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__10_ ( .D(aes_core_keymem_n2247), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[650]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__13_ ( .D(aes_core_keymem_n2211), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[653]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__14_ ( .D(aes_core_keymem_n2199), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[654]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__15_ ( .D(aes_core_keymem_n2187), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[655]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__16_ ( .D(aes_core_keymem_n2175), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[656]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__24_ ( .D(aes_core_keymem_n2079), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[664]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__26_ ( .D(aes_core_keymem_n2055), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[666]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__29_ ( .D(aes_core_keymem_n2019), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[669]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__30_ ( .D(aes_core_keymem_n2007), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[670]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__31_ ( .D(aes_core_keymem_n1995), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[671]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__32_ ( .D(aes_core_keymem_n1983), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[672]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__40_ ( .D(aes_core_keymem_n1887), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[680]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__42_ ( .D(aes_core_keymem_n1863), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[682]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__45_ ( .D(aes_core_keymem_n1827), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[685]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__46_ ( .D(aes_core_keymem_n1815), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[686]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__47_ ( .D(aes_core_keymem_n1803), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[687]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__48_ ( .D(aes_core_keymem_n1791), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[688]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__56_ ( .D(aes_core_keymem_n1695), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[696]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__58_ ( .D(aes_core_keymem_n1671), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[698]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__61_ ( .D(aes_core_keymem_n1635), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[701]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__62_ ( .D(aes_core_keymem_n1623), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[702]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__63_ ( .D(aes_core_keymem_n1611), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[703]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__64_ ( .D(aes_core_keymem_n1599), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[704]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__72_ ( .D(aes_core_keymem_n1503), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[712]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__74_ ( .D(aes_core_keymem_n1479), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[714]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__77_ ( .D(aes_core_keymem_n1443), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[717]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__78_ ( .D(aes_core_keymem_n1431), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[718]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__79_ ( .D(aes_core_keymem_n1419), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[719]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__80_ ( .D(aes_core_keymem_n1407), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[720]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__88_ ( .D(aes_core_keymem_n1311), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[728]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__90_ ( .D(aes_core_keymem_n1287), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[730]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__93_ ( .D(aes_core_keymem_n1251), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[733]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__94_ ( .D(aes_core_keymem_n1239), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[734]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__95_ ( .D(aes_core_keymem_n1227), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[735]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__96_ ( .D(aes_core_keymem_n1215), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[736]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__104_ ( .D(aes_core_keymem_n1119), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[744]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__106_ ( .D(aes_core_keymem_n1095), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[746]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__109_ ( .D(aes_core_keymem_n1059), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[749]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__110_ ( .D(aes_core_keymem_n1047), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[750]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__111_ ( .D(aes_core_keymem_n1035), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[751]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__112_ ( .D(aes_core_keymem_n1023), 
        .CK(clk_48Mhz), .Q(aes_core_keymem_key_mem[752]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__120_ ( .D(aes_core_keymem_n927), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[760]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__122_ ( .D(aes_core_keymem_n903), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[762]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__125_ ( .D(aes_core_keymem_n867), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[765]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__126_ ( .D(aes_core_keymem_n855), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[766]) );
  DFFHQX1 aes_core_keymem_key_mem_reg_9__127_ ( .D(aes_core_keymem_n843), .CK(
        clk_48Mhz), .Q(aes_core_keymem_key_mem[767]) );
  CLKINVX4 aes_core_keymem_U2519 ( .A(reset_n), .Y(aes_core_keymem_n14) );
  CLKINVX4 aes_core_keymem_U2515 ( .A(aes_core_keymem_n822), .Y(
        aes_core_keymem_n9) );
  NOR2X4 aes_core_keymem_U2465 ( .A(aes_core_keymem_n22), .B(
        aes_core_keymem_n14), .Y(aes_core_keymem_n822) );
  NAND4X4 aes_core_keymem_U2456 ( .A(aes_core_keymem_n826), .B(
        aes_core_keymem_n822), .C(aes_core_keymem_n2767), .D(
        aes_core_keymem_n2768), .Y(aes_core_keymem_n553) );
  NAND3X4 aes_core_keymem_U2454 ( .A(aes_core_keymem_n824), .B(
        aes_core_keymem_n822), .C(aes_core_keymem_n826), .Y(
        aes_core_keymem_n552) );
  NAND3X4 aes_core_keymem_U2452 ( .A(aes_core_keymem_n822), .B(
        aes_core_keymem_n827), .C(aes_core_keymem_n826), .Y(
        aes_core_keymem_n551) );
  NAND3X4 aes_core_keymem_U2450 ( .A(aes_core_keymem_n825), .B(
        aes_core_keymem_n822), .C(aes_core_keymem_n826), .Y(
        aes_core_keymem_n550) );
  NAND4X4 aes_core_keymem_U2448 ( .A(aes_core_keymem_n822), .B(
        aes_core_keymem_n823), .C(aes_core_keymem_n2767), .D(
        aes_core_keymem_n2768), .Y(aes_core_keymem_n549) );
  NAND3X4 aes_core_keymem_U2446 ( .A(aes_core_keymem_n822), .B(
        aes_core_keymem_n823), .C(aes_core_keymem_n824), .Y(
        aes_core_keymem_n548) );
  OR2X4 aes_core_keymem_U2444 ( .A(aes_core_keymem_n821), .B(
        aes_core_keymem_n9), .Y(aes_core_keymem_n547) );
  DFFRHQX4 aes_core_keymem_key_mem_ctrl_reg_reg_1_ ( .D(aes_core_keymem_n2388), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem_ctrl_reg[1])
         );
  DFFRHQX4 aes_core_keymem_key_mem_ctrl_reg_reg_0_ ( .D(aes_core_keymem_n2390), 
        .CK(clk_48Mhz), .RN(reset_n), .Q(aes_core_keymem_key_mem_ctrl_reg[0])
         );
  BUFX3 aes_core_sbox_inst_U1767 ( .A(aes_core_n24), .Y(aes_core_sbox_inst_n62) );
  BUFX3 aes_core_sbox_inst_U1766 ( .A(aes_core_n8), .Y(aes_core_sbox_inst_n56)
         );
  BUFX3 aes_core_sbox_inst_U1765 ( .A(aes_core_n32), .Y(aes_core_sbox_inst_n64) );
  BUFX3 aes_core_sbox_inst_U1764 ( .A(aes_core_n28), .Y(aes_core_sbox_inst_n63) );
  NOR2X1 aes_core_sbox_inst_U1763 ( .A(aes_core_sbox_inst_n206), .B(
        aes_core_sbox_inst_n64), .Y(aes_core_sbox_inst_n839) );
  NOR2X1 aes_core_sbox_inst_U1762 ( .A(aes_core_sbox_inst_n148), .B(
        aes_core_sbox_inst_n64), .Y(aes_core_sbox_inst_n673) );
  NOR2X1 aes_core_sbox_inst_U1761 ( .A(aes_core_sbox_inst_n58), .B(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n271) );
  BUFX3 aes_core_sbox_inst_U1760 ( .A(aes_core_sbox_inst_n271), .Y(
        aes_core_sbox_inst_n84) );
  NAND2X1 aes_core_sbox_inst_U1759 ( .A(aes_core_sbox_inst_n315), .B(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n1391) );
  NOR2X1 aes_core_sbox_inst_U1758 ( .A(aes_core_sbox_inst_n1682), .B(
        aes_core_sbox_inst_n56), .Y(aes_core_sbox_inst_n572) );
  NOR2X1 aes_core_sbox_inst_U1757 ( .A(aes_core_sbox_inst_n450), .B(
        aes_core_sbox_inst_n62), .Y(aes_core_sbox_inst_n1197) );
  NOR2X1 aes_core_sbox_inst_U1756 ( .A(aes_core_sbox_inst_n1620), .B(
        aes_core_n16), .Y(aes_core_sbox_inst_n1478) );
  NOR2X1 aes_core_sbox_inst_U1755 ( .A(aes_core_sbox_inst_n59), .B(
        aes_core_n14), .Y(aes_core_sbox_inst_n275) );
  OAI22X1 aes_core_sbox_inst_U1754 ( .A0(aes_core_sbox_inst_n38), .A1(
        aes_core_sbox_inst_n42), .B0(aes_core_sbox_inst_n58), .B1(
        aes_core_sbox_inst_n33), .Y(aes_core_sbox_inst_n294) );
  NOR2X1 aes_core_sbox_inst_U1753 ( .A(aes_core_sbox_inst_n34), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n345) );
  OAI221X1 aes_core_sbox_inst_U1752 ( .A0(aes_core_sbox_inst_n107), .A1(
        aes_core_sbox_inst_n15), .B0(aes_core_n30), .B1(
        aes_core_sbox_inst_n160), .C0(aes_core_n29), .Y(
        aes_core_sbox_inst_n763) );
  OAI221X1 aes_core_sbox_inst_U1751 ( .A0(aes_core_sbox_inst_n79), .A1(
        aes_core_sbox_inst_n34), .B0(aes_core_sbox_inst_n57), .B1(aes_core_n14), .C0(aes_core_n13), .Y(aes_core_sbox_inst_n1411) );
  NOR2X1 aes_core_sbox_inst_U1750 ( .A(aes_core_sbox_inst_n39), .B(
        aes_core_n14), .Y(aes_core_sbox_inst_n367) );
  NOR2X1 aes_core_sbox_inst_U1749 ( .A(aes_core_sbox_inst_n51), .B(aes_core_n6), .Y(aes_core_sbox_inst_n545) );
  NOR2X1 aes_core_sbox_inst_U1748 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_sbox_inst_n61), .Y(aes_core_sbox_inst_n1140) );
  NOR2X1 aes_core_sbox_inst_U1747 ( .A(aes_core_sbox_inst_n18), .B(
        aes_core_n30), .Y(aes_core_sbox_inst_n812) );
  NOR2X1 aes_core_sbox_inst_U1746 ( .A(aes_core_sbox_inst_n59), .B(
        aes_core_n13), .Y(aes_core_sbox_inst_n314) );
  NOR2X1 aes_core_sbox_inst_U1745 ( .A(aes_core_sbox_inst_n55), .B(aes_core_n5), .Y(aes_core_sbox_inst_n410) );
  NOR2X1 aes_core_sbox_inst_U1744 ( .A(aes_core_sbox_inst_n60), .B(
        aes_core_n21), .Y(aes_core_sbox_inst_n1005) );
  NOR2X1 aes_core_sbox_inst_U1743 ( .A(aes_core_sbox_inst_n63), .B(
        aes_core_n29), .Y(aes_core_sbox_inst_n643) );
  NOR2X1 aes_core_sbox_inst_U1742 ( .A(aes_core_sbox_inst_n186), .B(
        aes_core_sbox_inst_n56), .Y(aes_core_sbox_inst_n529) );
  NOR2X1 aes_core_sbox_inst_U1741 ( .A(aes_core_sbox_inst_n164), .B(
        aes_core_sbox_inst_n62), .Y(aes_core_sbox_inst_n1124) );
  NOR2X1 aes_core_sbox_inst_U1740 ( .A(aes_core_sbox_inst_n146), .B(
        aes_core_sbox_inst_n64), .Y(aes_core_sbox_inst_n796) );
  NOR2X1 aes_core_sbox_inst_U1739 ( .A(aes_core_sbox_inst_n179), .B(
        aes_core_n16), .Y(aes_core_sbox_inst_n1372) );
  NOR2X1 aes_core_sbox_inst_U1738 ( .A(aes_core_sbox_inst_n166), .B(
        aes_core_sbox_inst_n62), .Y(aes_core_sbox_inst_n1035) );
  INVX1 aes_core_sbox_inst_U1737 ( .A(aes_core_n7), .Y(aes_core_sbox_inst_n189) );
  NAND3X1 aes_core_sbox_inst_U1736 ( .A(aes_core_sbox_inst_n1704), .B(
        aes_core_sbox_inst_n126), .C(aes_core_sbox_inst_n55), .Y(
        aes_core_sbox_inst_n554) );
  NAND3X1 aes_core_sbox_inst_U1735 ( .A(aes_core_sbox_inst_n1586), .B(
        aes_core_sbox_inst_n121), .C(aes_core_sbox_inst_n60), .Y(
        aes_core_sbox_inst_n1149) );
  NAND4X1 aes_core_sbox_inst_U1734 ( .A(aes_core_sbox_inst_n1148), .B(
        aes_core_sbox_inst_n990), .C(aes_core_sbox_inst_n1149), .D(
        aes_core_sbox_inst_n1150), .Y(aes_core_sbox_inst_n1147) );
  AOI22X1 aes_core_sbox_inst_U1733 ( .A0(aes_core_sbox_inst_n1048), .A1(
        aes_core_sbox_inst_n4), .B0(aes_core_sbox_inst_n1124), .B1(
        aes_core_sbox_inst_n1147), .Y(aes_core_sbox_inst_n1146) );
  INVX1 aes_core_sbox_inst_U1732 ( .A(aes_core_sbox_inst_n1146), .Y(
        aes_core_sbox_inst_n1570) );
  NAND3X1 aes_core_sbox_inst_U1731 ( .A(aes_core_sbox_inst_n227), .B(
        aes_core_sbox_inst_n117), .C(aes_core_sbox_inst_n63), .Y(
        aes_core_sbox_inst_n821) );
  NAND4X1 aes_core_sbox_inst_U1730 ( .A(aes_core_sbox_inst_n820), .B(
        aes_core_sbox_inst_n628), .C(aes_core_sbox_inst_n821), .D(
        aes_core_sbox_inst_n822), .Y(aes_core_sbox_inst_n819) );
  AOI22X1 aes_core_sbox_inst_U1729 ( .A0(aes_core_sbox_inst_n686), .A1(
        aes_core_sbox_inst_n9), .B0(aes_core_sbox_inst_n796), .B1(
        aes_core_sbox_inst_n819), .Y(aes_core_sbox_inst_n818) );
  INVX1 aes_core_sbox_inst_U1728 ( .A(aes_core_sbox_inst_n818), .Y(
        aes_core_sbox_inst_n212) );
  XNOR2X1 aes_core_sbox_inst_U1727 ( .A(aes_core_sbox_inst_n55), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n1563) );
  NAND2X1 aes_core_sbox_inst_U1726 ( .A(aes_core_sbox_inst_n1563), .B(
        aes_core_sbox_inst_n1735), .Y(aes_core_sbox_inst_n1545) );
  XNOR2X1 aes_core_sbox_inst_U1725 ( .A(aes_core_sbox_inst_n60), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1321) );
  NAND2X1 aes_core_sbox_inst_U1724 ( .A(aes_core_sbox_inst_n1321), .B(
        aes_core_sbox_inst_n30), .Y(aes_core_sbox_inst_n1303) );
  XNOR2X1 aes_core_sbox_inst_U1723 ( .A(aes_core_sbox_inst_n63), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n963) );
  NAND2X1 aes_core_sbox_inst_U1722 ( .A(aes_core_sbox_inst_n963), .B(
        aes_core_sbox_inst_n20), .Y(aes_core_sbox_inst_n945) );
  AOI222X1 aes_core_sbox_inst_U1721 ( .A0(aes_core_sbox_inst_n77), .A1(
        aes_core_sbox_inst_n128), .B0(aes_core_sbox_inst_n538), .B1(
        aes_core_sbox_inst_n192), .C0(aes_core_sbox_inst_n76), .C1(
        aes_core_sbox_inst_n67), .Y(aes_core_sbox_inst_n537) );
  NAND3X1 aes_core_sbox_inst_U1720 ( .A(aes_core_sbox_inst_n55), .B(
        aes_core_sbox_inst_n126), .C(aes_core_sbox_inst_n385), .Y(
        aes_core_sbox_inst_n536) );
  NAND4X1 aes_core_sbox_inst_U1719 ( .A(aes_core_sbox_inst_n534), .B(
        aes_core_sbox_inst_n535), .C(aes_core_sbox_inst_n536), .D(
        aes_core_sbox_inst_n537), .Y(aes_core_sbox_inst_n530) );
  AOI222X1 aes_core_sbox_inst_U1718 ( .A0(aes_core_sbox_inst_n103), .A1(
        aes_core_sbox_inst_n123), .B0(aes_core_sbox_inst_n1133), .B1(
        aes_core_sbox_inst_n170), .C0(aes_core_sbox_inst_n102), .C1(
        aes_core_sbox_inst_n93), .Y(aes_core_sbox_inst_n1132) );
  NAND3X1 aes_core_sbox_inst_U1717 ( .A(aes_core_sbox_inst_n60), .B(
        aes_core_sbox_inst_n121), .C(aes_core_sbox_inst_n980), .Y(
        aes_core_sbox_inst_n1131) );
  NAND4X1 aes_core_sbox_inst_U1716 ( .A(aes_core_sbox_inst_n1129), .B(
        aes_core_sbox_inst_n1130), .C(aes_core_sbox_inst_n1131), .D(
        aes_core_sbox_inst_n1132), .Y(aes_core_sbox_inst_n1125) );
  AOI222X1 aes_core_sbox_inst_U1715 ( .A0(aes_core_sbox_inst_n115), .A1(
        aes_core_sbox_inst_n119), .B0(aes_core_sbox_inst_n805), .B1(
        aes_core_sbox_inst_n154), .C0(aes_core_sbox_inst_n114), .C1(
        aes_core_sbox_inst_n107), .Y(aes_core_sbox_inst_n804) );
  NAND3X1 aes_core_sbox_inst_U1714 ( .A(aes_core_sbox_inst_n63), .B(
        aes_core_sbox_inst_n117), .C(aes_core_sbox_inst_n618), .Y(
        aes_core_sbox_inst_n803) );
  NAND4X1 aes_core_sbox_inst_U1713 ( .A(aes_core_sbox_inst_n801), .B(
        aes_core_sbox_inst_n802), .C(aes_core_sbox_inst_n803), .D(
        aes_core_sbox_inst_n804), .Y(aes_core_sbox_inst_n797) );
  AOI222X1 aes_core_sbox_inst_U1712 ( .A0(aes_core_sbox_inst_n57), .A1(
        aes_core_sbox_inst_n85), .B0(aes_core_sbox_inst_n367), .B1(
        aes_core_sbox_inst_n79), .C0(aes_core_sbox_inst_n143), .C1(
        aes_core_sbox_inst_n90), .Y(aes_core_sbox_inst_n366) );
  AOI21X1 aes_core_sbox_inst_U1711 ( .A0(aes_core_sbox_inst_n368), .A1(
        aes_core_sbox_inst_n1656), .B0(aes_core_sbox_inst_n369), .Y(
        aes_core_sbox_inst_n365) );
  NAND4X1 aes_core_sbox_inst_U1710 ( .A(aes_core_sbox_inst_n320), .B(
        aes_core_sbox_inst_n36), .C(aes_core_sbox_inst_n365), .D(
        aes_core_sbox_inst_n366), .Y(aes_core_sbox_inst_n363) );
  AOI222X1 aes_core_sbox_inst_U1709 ( .A0(aes_core_sbox_inst_n83), .A1(
        aes_core_sbox_inst_n45), .B0(aes_core_sbox_inst_n276), .B1(
        aes_core_sbox_inst_n58), .C0(aes_core_sbox_inst_n89), .C1(
        aes_core_sbox_inst_n79), .Y(aes_core_sbox_inst_n1449) );
  NAND3X1 aes_core_sbox_inst_U1708 ( .A(aes_core_sbox_inst_n59), .B(
        aes_core_sbox_inst_n41), .C(aes_core_sbox_inst_n1446), .Y(
        aes_core_sbox_inst_n1448) );
  NAND4X1 aes_core_sbox_inst_U1707 ( .A(aes_core_sbox_inst_n1447), .B(
        aes_core_sbox_inst_n319), .C(aes_core_sbox_inst_n1448), .D(
        aes_core_sbox_inst_n1449), .Y(aes_core_sbox_inst_n1442) );
  AOI22X1 aes_core_sbox_inst_U1706 ( .A0(aes_core_sbox_inst_n283), .A1(
        aes_core_sbox_inst_n1678), .B0(aes_core_sbox_inst_n57), .B1(
        aes_core_sbox_inst_n272), .Y(aes_core_sbox_inst_n278) );
  AOI222X1 aes_core_sbox_inst_U1705 ( .A0(aes_core_sbox_inst_n88), .A1(
        aes_core_sbox_inst_n84), .B0(aes_core_sbox_inst_n90), .B1(
        aes_core_sbox_inst_n125), .C0(aes_core_sbox_inst_n79), .C1(
        aes_core_sbox_inst_n83), .Y(aes_core_sbox_inst_n279) );
  NAND4BX1 aes_core_sbox_inst_U1704 ( .AN(aes_core_sbox_inst_n277), .B(
        aes_core_sbox_inst_n1666), .C(aes_core_sbox_inst_n278), .D(
        aes_core_sbox_inst_n279), .Y(aes_core_sbox_inst_n264) );
  NOR2X1 aes_core_sbox_inst_U1703 ( .A(aes_core_sbox_inst_n1720), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n382) );
  BUFX3 aes_core_sbox_inst_U1702 ( .A(aes_core_sbox_inst_n382), .Y(
        aes_core_sbox_inst_n76) );
  AOI222X1 aes_core_sbox_inst_U1701 ( .A0(aes_core_sbox_inst_n82), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n84), .B1(
        aes_core_sbox_inst_n272), .C0(aes_core_sbox_inst_n143), .C1(
        aes_core_sbox_inst_n88), .Y(aes_core_sbox_inst_n269) );
  AOI22X1 aes_core_sbox_inst_U1700 ( .A0(aes_core_sbox_inst_n275), .A1(
        aes_core_sbox_inst_n57), .B0(aes_core_sbox_inst_n276), .B1(
        aes_core_sbox_inst_n144), .Y(aes_core_sbox_inst_n268) );
  NAND4BX1 aes_core_sbox_inst_U1699 ( .AN(aes_core_sbox_inst_n267), .B(
        aes_core_sbox_inst_n1668), .C(aes_core_sbox_inst_n268), .D(
        aes_core_sbox_inst_n269), .Y(aes_core_sbox_inst_n266) );
  NOR2X1 aes_core_sbox_inst_U1698 ( .A(aes_core_sbox_inst_n24), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n977) );
  BUFX3 aes_core_sbox_inst_U1697 ( .A(aes_core_sbox_inst_n977), .Y(
        aes_core_sbox_inst_n102) );
  INVX1 aes_core_sbox_inst_U1696 ( .A(aes_core_sbox_inst_n12), .Y(
        aes_core_sbox_inst_n1045) );
  OR2X2 aes_core_sbox_inst_U1695 ( .A(aes_core_sbox_inst_n22), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n12) );
  NOR2X1 aes_core_sbox_inst_U1694 ( .A(aes_core_sbox_inst_n243), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n615) );
  BUFX3 aes_core_sbox_inst_U1693 ( .A(aes_core_sbox_inst_n615), .Y(
        aes_core_sbox_inst_n114) );
  INVX1 aes_core_sbox_inst_U1692 ( .A(aes_core_sbox_inst_n11), .Y(
        aes_core_sbox_inst_n683) );
  OR2X2 aes_core_sbox_inst_U1691 ( .A(aes_core_sbox_inst_n14), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n11) );
  NOR2X1 aes_core_sbox_inst_U1690 ( .A(aes_core_sbox_inst_n37), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n357) );
  BUFX3 aes_core_sbox_inst_U1689 ( .A(aes_core_sbox_inst_n357), .Y(
        aes_core_sbox_inst_n89) );
  AOI22X1 aes_core_sbox_inst_U1688 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n57), .B0(aes_core_sbox_inst_n81), .B1(
        aes_core_sbox_inst_n90), .Y(aes_core_sbox_inst_n1489) );
  AOI22X1 aes_core_sbox_inst_U1687 ( .A0(aes_core_sbox_inst_n344), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n313), .B1(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n1525) );
  NOR2X1 aes_core_sbox_inst_U1686 ( .A(aes_core_n29), .B(aes_core_n30), .Y(
        aes_core_sbox_inst_n712) );
  BUFX3 aes_core_sbox_inst_U1685 ( .A(aes_core_sbox_inst_n712), .Y(
        aes_core_sbox_inst_n110) );
  NOR2X1 aes_core_sbox_inst_U1684 ( .A(aes_core_sbox_inst_n127), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n448) );
  NOR2X1 aes_core_sbox_inst_U1683 ( .A(aes_core_sbox_inst_n122), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1043) );
  NOR2X1 aes_core_sbox_inst_U1682 ( .A(aes_core_sbox_inst_n118), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n681) );
  AOI22X1 aes_core_sbox_inst_U1681 ( .A0(aes_core_sbox_inst_n276), .A1(
        aes_core_sbox_inst_n44), .B0(aes_core_sbox_inst_n83), .B1(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n341) );
  AOI31X1 aes_core_sbox_inst_U1680 ( .A0(aes_core_sbox_inst_n341), .A1(
        aes_core_sbox_inst_n342), .A2(aes_core_sbox_inst_n343), .B0(
        aes_core_sbox_inst_n181), .Y(aes_core_sbox_inst_n339) );
  NOR3X1 aes_core_sbox_inst_U1679 ( .A(aes_core_sbox_inst_n31), .B(
        aes_core_n13), .C(aes_core_sbox_inst_n40), .Y(aes_core_sbox_inst_n340)
         );
  NOR3BX1 aes_core_sbox_inst_U1678 ( .AN(aes_core_sbox_inst_n338), .B(
        aes_core_sbox_inst_n339), .C(aes_core_sbox_inst_n340), .Y(
        aes_core_sbox_inst_n325) );
  AOI22X1 aes_core_sbox_inst_U1677 ( .A0(aes_core_sbox_inst_n561), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n508), .B1(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n749) );
  AOI22X1 aes_core_sbox_inst_U1676 ( .A0(aes_core_sbox_inst_n1156), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n1103), .B1(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1254) );
  AOI22X1 aes_core_sbox_inst_U1675 ( .A0(aes_core_sbox_inst_n828), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n775), .B1(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n896) );
  NOR2X1 aes_core_sbox_inst_U1674 ( .A(aes_core_sbox_inst_n35), .B(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n1363) );
  NAND2X1 aes_core_sbox_inst_U1673 ( .A(aes_core_sbox_inst_n83), .B(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n1348) );
  NAND3X1 aes_core_sbox_inst_U1672 ( .A(aes_core_n6), .B(
        aes_core_sbox_inst_n1732), .C(aes_core_sbox_inst_n139), .Y(
        aes_core_sbox_inst_n534) );
  NAND3X1 aes_core_sbox_inst_U1671 ( .A(aes_core_sbox_inst_n61), .B(
        aes_core_sbox_inst_n27), .C(aes_core_sbox_inst_n130), .Y(
        aes_core_sbox_inst_n1129) );
  NAND3X1 aes_core_sbox_inst_U1670 ( .A(aes_core_n30), .B(
        aes_core_sbox_inst_n18), .C(aes_core_sbox_inst_n135), .Y(
        aes_core_sbox_inst_n801) );
  AOI31X1 aes_core_sbox_inst_U1669 ( .A0(aes_core_sbox_inst_n139), .A1(
        aes_core_n6), .A2(aes_core_sbox_inst_n399), .B0(
        aes_core_sbox_inst_n464), .Y(aes_core_sbox_inst_n1559) );
  AOI31X1 aes_core_sbox_inst_U1668 ( .A0(aes_core_sbox_inst_n130), .A1(
        aes_core_sbox_inst_n61), .A2(aes_core_sbox_inst_n994), .B0(
        aes_core_sbox_inst_n1059), .Y(aes_core_sbox_inst_n1317) );
  AOI31X1 aes_core_sbox_inst_U1667 ( .A0(aes_core_sbox_inst_n135), .A1(
        aes_core_n30), .A2(aes_core_sbox_inst_n632), .B0(
        aes_core_sbox_inst_n697), .Y(aes_core_sbox_inst_n959) );
  AOI22X1 aes_core_sbox_inst_U1666 ( .A0(aes_core_sbox_inst_n51), .A1(
        aes_core_sbox_inst_n201), .B0(aes_core_sbox_inst_n55), .B1(
        aes_core_sbox_inst_n5), .Y(aes_core_sbox_inst_n580) );
  AOI22X1 aes_core_sbox_inst_U1665 ( .A0(aes_core_sbox_inst_n26), .A1(
        aes_core_sbox_inst_n175), .B0(aes_core_sbox_inst_n60), .B1(
        aes_core_sbox_inst_n4), .Y(aes_core_sbox_inst_n1205) );
  AOI22X1 aes_core_sbox_inst_U1664 ( .A0(aes_core_sbox_inst_n18), .A1(
        aes_core_sbox_inst_n161), .B0(aes_core_sbox_inst_n63), .B1(
        aes_core_sbox_inst_n9), .Y(aes_core_sbox_inst_n847) );
  AOI22X1 aes_core_sbox_inst_U1663 ( .A0(aes_core_sbox_inst_n39), .A1(
        aes_core_sbox_inst_n57), .B0(aes_core_sbox_inst_n2), .B1(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n336) );
  AOI22X1 aes_core_sbox_inst_U1662 ( .A0(aes_core_sbox_inst_n86), .A1(
        aes_core_sbox_inst_n58), .B0(aes_core_sbox_inst_n40), .B1(
        aes_core_sbox_inst_n83), .Y(aes_core_sbox_inst_n1514) );
  INVX1 aes_core_sbox_inst_U1661 ( .A(aes_core_sbox_inst_n581), .Y(
        aes_core_sbox_inst_n1689) );
  AOI31X1 aes_core_sbox_inst_U1660 ( .A0(aes_core_sbox_inst_n199), .A1(
        aes_core_n6), .A2(aes_core_sbox_inst_n399), .B0(
        aes_core_sbox_inst_n1689), .Y(aes_core_sbox_inst_n569) );
  INVX1 aes_core_sbox_inst_U1659 ( .A(aes_core_sbox_inst_n1206), .Y(
        aes_core_sbox_inst_n1571) );
  AOI31X1 aes_core_sbox_inst_U1658 ( .A0(aes_core_sbox_inst_n174), .A1(
        aes_core_sbox_inst_n61), .A2(aes_core_sbox_inst_n994), .B0(
        aes_core_sbox_inst_n1571), .Y(aes_core_sbox_inst_n1194) );
  INVX1 aes_core_sbox_inst_U1657 ( .A(aes_core_sbox_inst_n848), .Y(
        aes_core_sbox_inst_n213) );
  AOI31X1 aes_core_sbox_inst_U1656 ( .A0(aes_core_sbox_inst_n159), .A1(
        aes_core_n30), .A2(aes_core_sbox_inst_n632), .B0(
        aes_core_sbox_inst_n213), .Y(aes_core_sbox_inst_n836) );
  AOI22X1 aes_core_sbox_inst_U1655 ( .A0(aes_core_sbox_inst_n191), .A1(
        aes_core_sbox_inst_n55), .B0(aes_core_sbox_inst_n51), .B1(
        aes_core_sbox_inst_n383), .Y(aes_core_sbox_inst_n490) );
  AOI22X1 aes_core_sbox_inst_U1654 ( .A0(aes_core_sbox_inst_n169), .A1(
        aes_core_sbox_inst_n60), .B0(aes_core_sbox_inst_n26), .B1(
        aes_core_sbox_inst_n978), .Y(aes_core_sbox_inst_n1085) );
  AOI22X1 aes_core_sbox_inst_U1653 ( .A0(aes_core_sbox_inst_n151), .A1(
        aes_core_sbox_inst_n63), .B0(aes_core_sbox_inst_n18), .B1(
        aes_core_sbox_inst_n616), .Y(aes_core_sbox_inst_n723) );
  AOI22X1 aes_core_sbox_inst_U1652 ( .A0(aes_core_sbox_inst_n46), .A1(
        aes_core_sbox_inst_n39), .B0(aes_core_sbox_inst_n59), .B1(
        aes_core_sbox_inst_n80), .Y(aes_core_sbox_inst_n1393) );
  NOR2X1 aes_core_sbox_inst_U1651 ( .A(aes_core_sbox_inst_n150), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n721) );
  NOR2X1 aes_core_sbox_inst_U1650 ( .A(aes_core_sbox_inst_n67), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n463) );
  NOR2X1 aes_core_sbox_inst_U1649 ( .A(aes_core_sbox_inst_n93), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1058) );
  NOR2X1 aes_core_sbox_inst_U1648 ( .A(aes_core_sbox_inst_n107), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n696) );
  NOR2X1 aes_core_sbox_inst_U1647 ( .A(aes_core_sbox_inst_n79), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n368) );
  OAI221X1 aes_core_sbox_inst_U1646 ( .A0(aes_core_sbox_inst_n67), .A1(
        aes_core_sbox_inst_n49), .B0(aes_core_n6), .B1(aes_core_sbox_inst_n196), .C0(aes_core_n5), .Y(aes_core_sbox_inst_n496) );
  OAI221X1 aes_core_sbox_inst_U1645 ( .A0(aes_core_sbox_inst_n93), .A1(
        aes_core_sbox_inst_n23), .B0(aes_core_sbox_inst_n61), .B1(
        aes_core_sbox_inst_n174), .C0(aes_core_n21), .Y(
        aes_core_sbox_inst_n1091) );
  OAI22X1 aes_core_sbox_inst_U1644 ( .A0(aes_core_sbox_inst_n59), .A1(
        aes_core_sbox_inst_n80), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n296) );
  OAI22X1 aes_core_sbox_inst_U1643 ( .A0(aes_core_sbox_inst_n138), .A1(
        aes_core_sbox_inst_n51), .B0(aes_core_sbox_inst_n55), .B1(
        aes_core_sbox_inst_n6), .Y(aes_core_sbox_inst_n406) );
  OAI22X1 aes_core_sbox_inst_U1642 ( .A0(aes_core_sbox_inst_n129), .A1(
        aes_core_sbox_inst_n26), .B0(aes_core_sbox_inst_n60), .B1(
        aes_core_sbox_inst_n7), .Y(aes_core_sbox_inst_n1001) );
  OAI22X1 aes_core_sbox_inst_U1641 ( .A0(aes_core_sbox_inst_n134), .A1(
        aes_core_sbox_inst_n18), .B0(aes_core_sbox_inst_n63), .B1(
        aes_core_sbox_inst_n8), .Y(aes_core_sbox_inst_n639) );
  AOI222X1 aes_core_sbox_inst_U1640 ( .A0(aes_core_sbox_inst_n313), .A1(
        aes_core_sbox_inst_n59), .B0(aes_core_sbox_inst_n314), .B1(
        aes_core_sbox_inst_n79), .C0(aes_core_sbox_inst_n315), .C1(
        aes_core_sbox_inst_n43), .Y(aes_core_sbox_inst_n312) );
  AOI222X1 aes_core_sbox_inst_U1639 ( .A0(aes_core_sbox_inst_n84), .A1(
        aes_core_sbox_inst_n321), .B0(aes_core_sbox_inst_n344), .B1(
        aes_core_sbox_inst_n79), .C0(aes_core_sbox_inst_n57), .C1(
        aes_core_sbox_inst_n10), .Y(aes_core_sbox_inst_n1468) );
  NOR2X1 aes_core_sbox_inst_U1638 ( .A(aes_core_sbox_inst_n50), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n538) );
  NOR2X1 aes_core_sbox_inst_U1637 ( .A(aes_core_sbox_inst_n25), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1133) );
  NOR2X1 aes_core_sbox_inst_U1636 ( .A(aes_core_sbox_inst_n17), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n805) );
  AOI211X1 aes_core_sbox_inst_U1635 ( .A0(aes_core_sbox_inst_n1379), .A1(
        aes_core_sbox_inst_n58), .B0(aes_core_sbox_inst_n83), .C0(
        aes_core_sbox_inst_n1356), .Y(aes_core_sbox_inst_n1460) );
  AOI222X1 aes_core_sbox_inst_U1634 ( .A0(aes_core_sbox_inst_n88), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n57), .B1(
        aes_core_sbox_inst_n10), .C0(aes_core_sbox_inst_n90), .C1(
        aes_core_sbox_inst_n47), .Y(aes_core_sbox_inst_n1497) );
  AOI222X1 aes_core_sbox_inst_U1633 ( .A0(aes_core_sbox_inst_n508), .A1(
        aes_core_sbox_inst_n55), .B0(aes_core_sbox_inst_n410), .B1(
        aes_core_sbox_inst_n67), .C0(aes_core_sbox_inst_n469), .C1(
        aes_core_sbox_inst_n193), .Y(aes_core_sbox_inst_n1188) );
  AOI222X1 aes_core_sbox_inst_U1632 ( .A0(aes_core_sbox_inst_n1103), .A1(
        aes_core_sbox_inst_n60), .B0(aes_core_sbox_inst_n1005), .B1(
        aes_core_sbox_inst_n93), .C0(aes_core_sbox_inst_n1064), .C1(
        aes_core_sbox_inst_n173), .Y(aes_core_sbox_inst_n1292) );
  AOI222X1 aes_core_sbox_inst_U1631 ( .A0(aes_core_sbox_inst_n775), .A1(
        aes_core_sbox_inst_n63), .B0(aes_core_sbox_inst_n643), .B1(
        aes_core_sbox_inst_n107), .C0(aes_core_sbox_inst_n702), .C1(
        aes_core_sbox_inst_n155), .Y(aes_core_sbox_inst_n934) );
  AOI22X1 aes_core_sbox_inst_U1630 ( .A0(aes_core_sbox_inst_n59), .A1(
        aes_core_sbox_inst_n58), .B0(aes_core_sbox_inst_n39), .B1(
        aes_core_sbox_inst_n80), .Y(aes_core_sbox_inst_n1404) );
  NAND2X1 aes_core_sbox_inst_U1629 ( .A(aes_core_sbox_inst_n37), .B(
        aes_core_sbox_inst_n1637), .Y(aes_core_sbox_inst_n1513) );
  AOI222X1 aes_core_sbox_inst_U1628 ( .A0(aes_core_sbox_inst_n90), .A1(
        aes_core_sbox_inst_n125), .B0(aes_core_sbox_inst_n58), .B1(
        aes_core_sbox_inst_n1513), .C0(aes_core_sbox_inst_n367), .C1(
        aes_core_sbox_inst_n80), .Y(aes_core_sbox_inst_n1512) );
  NOR2X1 aes_core_sbox_inst_U1627 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_n21), .Y(aes_core_sbox_inst_n1156) );
  NOR2X1 aes_core_sbox_inst_U1626 ( .A(aes_core_sbox_inst_n255), .B(
        aes_core_n29), .Y(aes_core_sbox_inst_n828) );
  INVX1 aes_core_sbox_inst_U1625 ( .A(aes_core_n15), .Y(
        aes_core_sbox_inst_n185) );
  INVX1 aes_core_sbox_inst_U1624 ( .A(aes_core_sbox_inst_n185), .Y(
        aes_core_sbox_inst_n183) );
  INVX1 aes_core_sbox_inst_U1623 ( .A(aes_core_n14), .Y(
        aes_core_sbox_inst_n1657) );
  BUFX3 aes_core_sbox_inst_U1622 ( .A(aes_core_sbox_inst_n1657), .Y(
        aes_core_sbox_inst_n34) );
  NAND3X1 aes_core_sbox_inst_U1621 ( .A(aes_core_sbox_inst_n1656), .B(
        aes_core_sbox_inst_n41), .C(aes_core_sbox_inst_n59), .Y(
        aes_core_sbox_inst_n1463) );
  INVX1 aes_core_sbox_inst_U1620 ( .A(aes_core_n30), .Y(
        aes_core_sbox_inst_n236) );
  INVX1 aes_core_sbox_inst_U1619 ( .A(aes_core_sbox_inst_n57), .Y(
        aes_core_sbox_inst_n1679) );
  INVX1 aes_core_sbox_inst_U1618 ( .A(aes_core_sbox_inst_n58), .Y(
        aes_core_sbox_inst_n1676) );
  INVX1 aes_core_sbox_inst_U1617 ( .A(aes_core_sbox_inst_n55), .Y(
        aes_core_sbox_inst_n1732) );
  INVX1 aes_core_sbox_inst_U1616 ( .A(aes_core_sbox_inst_n60), .Y(
        aes_core_sbox_inst_n1614) );
  INVX1 aes_core_sbox_inst_U1615 ( .A(aes_core_sbox_inst_n59), .Y(
        aes_core_sbox_inst_n1674) );
  NOR2X1 aes_core_sbox_inst_U1614 ( .A(aes_core_sbox_inst_n23), .B(
        aes_core_n21), .Y(aes_core_sbox_inst_n1102) );
  BUFX3 aes_core_sbox_inst_U1613 ( .A(aes_core_sbox_inst_n1102), .Y(
        aes_core_sbox_inst_n92) );
  NOR2X1 aes_core_sbox_inst_U1612 ( .A(aes_core_sbox_inst_n1607), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1029) );
  AND2X2 aes_core_sbox_inst_U1611 ( .A(aes_core_sbox_inst_n291), .B(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n1358) );
  NOR2X1 aes_core_sbox_inst_U1610 ( .A(aes_core_n21), .B(
        aes_core_sbox_inst_n61), .Y(aes_core_sbox_inst_n1074) );
  BUFX3 aes_core_sbox_inst_U1609 ( .A(aes_core_sbox_inst_n1074), .Y(
        aes_core_sbox_inst_n97) );
  AOI21X1 aes_core_sbox_inst_U1608 ( .A0(aes_core_sbox_inst_n36), .A1(
        aes_core_sbox_inst_n1638), .B0(aes_core_sbox_inst_n124), .Y(
        aes_core_sbox_inst_n1483) );
  AOI221X1 aes_core_sbox_inst_U1607 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n58), .B0(aes_core_sbox_inst_n275), .B1(
        aes_core_sbox_inst_n79), .C0(aes_core_sbox_inst_n1483), .Y(
        aes_core_sbox_inst_n1482) );
  AOI222X1 aes_core_sbox_inst_U1606 ( .A0(aes_core_sbox_inst_n1393), .A1(
        aes_core_sbox_inst_n321), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n83), .C0(aes_core_sbox_inst_n356), .C1(
        aes_core_sbox_inst_n45), .Y(aes_core_sbox_inst_n1481) );
  AOI21X1 aes_core_sbox_inst_U1605 ( .A0(aes_core_sbox_inst_n1481), .A1(
        aes_core_sbox_inst_n1482), .B0(aes_core_sbox_inst_n181), .Y(
        aes_core_sbox_inst_n1479) );
  AOI222X1 aes_core_sbox_inst_U1604 ( .A0(aes_core_sbox_inst_n356), .A1(
        aes_core_sbox_inst_n45), .B0(aes_core_sbox_inst_n314), .B1(
        aes_core_sbox_inst_n57), .C0(aes_core_sbox_inst_n90), .C1(
        aes_core_sbox_inst_n144), .Y(aes_core_sbox_inst_n1347) );
  NOR2BX1 aes_core_sbox_inst_U1603 ( .AN(aes_core_sbox_inst_n1348), .B(
        aes_core_sbox_inst_n89), .Y(aes_core_sbox_inst_n1346) );
  NAND4X1 aes_core_sbox_inst_U1602 ( .A(aes_core_sbox_inst_n296), .B(
        aes_core_sbox_inst_n1650), .C(aes_core_sbox_inst_n1346), .D(
        aes_core_sbox_inst_n1347), .Y(aes_core_sbox_inst_n1327) );
  NOR2X1 aes_core_sbox_inst_U1601 ( .A(aes_core_sbox_inst_n58), .B(
        aes_core_sbox_inst_n1628), .Y(aes_core_sbox_inst_n1351) );
  NOR2X1 aes_core_sbox_inst_U1600 ( .A(aes_core_sbox_inst_n25), .B(
        aes_core_sbox_inst_n61), .Y(aes_core_sbox_inst_n1015) );
  BUFX3 aes_core_sbox_inst_U1599 ( .A(aes_core_sbox_inst_n1015), .Y(
        aes_core_sbox_inst_n99) );
  NOR2X1 aes_core_sbox_inst_U1598 ( .A(aes_core_sbox_inst_n50), .B(aes_core_n6), .Y(aes_core_sbox_inst_n420) );
  BUFX3 aes_core_sbox_inst_U1597 ( .A(aes_core_sbox_inst_n420), .Y(
        aes_core_sbox_inst_n73) );
  NOR2X1 aes_core_sbox_inst_U1596 ( .A(aes_core_sbox_inst_n17), .B(
        aes_core_n30), .Y(aes_core_sbox_inst_n653) );
  BUFX3 aes_core_sbox_inst_U1595 ( .A(aes_core_sbox_inst_n653), .Y(
        aes_core_sbox_inst_n111) );
  OAI2BB1X1 aes_core_sbox_inst_U1594 ( .A0N(aes_core_sbox_inst_n54), .A1N(
        aes_core_n5), .B0(aes_core_sbox_inst_n137), .Y(aes_core_sbox_inst_n512) );
  OAI2BB1X1 aes_core_sbox_inst_U1593 ( .A0N(aes_core_sbox_inst_n30), .A1N(
        aes_core_n21), .B0(aes_core_sbox_inst_n131), .Y(
        aes_core_sbox_inst_n1107) );
  AOI211X1 aes_core_sbox_inst_U1592 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n1100), .C0(
        aes_core_sbox_inst_n1101), .Y(aes_core_sbox_inst_n1099) );
  AOI21X1 aes_core_sbox_inst_U1591 ( .A0(aes_core_sbox_inst_n999), .A1(
        aes_core_sbox_inst_n1107), .B0(aes_core_sbox_inst_n1018), .Y(
        aes_core_sbox_inst_n1098) );
  NAND4X1 aes_core_sbox_inst_U1590 ( .A(aes_core_sbox_inst_n1597), .B(
        aes_core_sbox_inst_n1097), .C(aes_core_sbox_inst_n1098), .D(
        aes_core_sbox_inst_n1099), .Y(aes_core_sbox_inst_n1096) );
  OAI2BB1X1 aes_core_sbox_inst_U1589 ( .A0N(aes_core_sbox_inst_n259), .A1N(
        aes_core_n29), .B0(aes_core_sbox_inst_n136), .Y(
        aes_core_sbox_inst_n779) );
  AOI211X1 aes_core_sbox_inst_U1588 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n772), .C0(
        aes_core_sbox_inst_n773), .Y(aes_core_sbox_inst_n771) );
  AOI21X1 aes_core_sbox_inst_U1587 ( .A0(aes_core_sbox_inst_n637), .A1(
        aes_core_sbox_inst_n779), .B0(aes_core_sbox_inst_n656), .Y(
        aes_core_sbox_inst_n770) );
  NAND4X1 aes_core_sbox_inst_U1586 ( .A(aes_core_sbox_inst_n238), .B(
        aes_core_sbox_inst_n769), .C(aes_core_sbox_inst_n770), .D(
        aes_core_sbox_inst_n771), .Y(aes_core_sbox_inst_n768) );
  NOR2X1 aes_core_sbox_inst_U1585 ( .A(aes_core_sbox_inst_n38), .B(
        aes_core_n14), .Y(aes_core_sbox_inst_n270) );
  BUFX3 aes_core_sbox_inst_U1584 ( .A(aes_core_sbox_inst_n270), .Y(
        aes_core_sbox_inst_n82) );
  AOI21X1 aes_core_sbox_inst_U1583 ( .A0(aes_core_n6), .A1(
        aes_core_sbox_inst_n404), .B0(aes_core_sbox_inst_n405), .Y(
        aes_core_sbox_inst_n403) );
  AOI21X1 aes_core_sbox_inst_U1582 ( .A0(aes_core_n30), .A1(
        aes_core_sbox_inst_n637), .B0(aes_core_sbox_inst_n638), .Y(
        aes_core_sbox_inst_n636) );
  NAND2X1 aes_core_sbox_inst_U1581 ( .A(aes_core_sbox_inst_n1397), .B(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n360) );
  NOR2X1 aes_core_sbox_inst_U1580 ( .A(aes_core_sbox_inst_n1725), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n434) );
  NOR2X1 aes_core_sbox_inst_U1579 ( .A(aes_core_sbox_inst_n248), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n667) );
  AOI21X1 aes_core_sbox_inst_U1578 ( .A0(aes_core_sbox_inst_n883), .A1(
        aes_core_sbox_inst_n884), .B0(aes_core_n33), .Y(
        aes_core_sbox_inst_n873) );
  NAND4X1 aes_core_sbox_inst_U1577 ( .A(aes_core_sbox_inst_n898), .B(
        aes_core_sbox_inst_n899), .C(aes_core_sbox_inst_n900), .D(
        aes_core_sbox_inst_n901), .Y(aes_core_sbox_inst_n872) );
  AOI211X1 aes_core_sbox_inst_U1576 ( .A0(aes_core_sbox_inst_n839), .A1(
        aes_core_sbox_inst_n872), .B0(aes_core_sbox_inst_n873), .C0(
        aes_core_sbox_inst_n874), .Y(aes_core_sbox_inst_n871) );
  INVX1 aes_core_sbox_inst_U1575 ( .A(aes_core_sbox_inst_n871), .Y(
        aes_core_new_sboxw[26]) );
  NOR2X1 aes_core_sbox_inst_U1574 ( .A(aes_core_n13), .B(aes_core_n14), .Y(
        aes_core_sbox_inst_n295) );
  BUFX3 aes_core_sbox_inst_U1573 ( .A(aes_core_sbox_inst_n295), .Y(
        aes_core_sbox_inst_n85) );
  NOR2X1 aes_core_sbox_inst_U1572 ( .A(aes_core_sbox_inst_n1645), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n280) );
  BUFX3 aes_core_sbox_inst_U1571 ( .A(aes_core_sbox_inst_n280), .Y(
        aes_core_sbox_inst_n90) );
  NOR2X1 aes_core_sbox_inst_U1570 ( .A(aes_core_sbox_inst_n1712), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n391) );
  BUFX3 aes_core_sbox_inst_U1569 ( .A(aes_core_sbox_inst_n391), .Y(
        aes_core_sbox_inst_n74) );
  NOR2X1 aes_core_sbox_inst_U1568 ( .A(aes_core_sbox_inst_n1594), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n986) );
  BUFX3 aes_core_sbox_inst_U1567 ( .A(aes_core_sbox_inst_n986), .Y(
        aes_core_sbox_inst_n100) );
  NOR2X1 aes_core_sbox_inst_U1566 ( .A(aes_core_sbox_inst_n235), .B(
        aes_core_sbox_inst_n63), .Y(aes_core_sbox_inst_n624) );
  BUFX3 aes_core_sbox_inst_U1565 ( .A(aes_core_sbox_inst_n624), .Y(
        aes_core_sbox_inst_n112) );
  NOR2X1 aes_core_sbox_inst_U1564 ( .A(aes_core_sbox_inst_n49), .B(aes_core_n5), .Y(aes_core_sbox_inst_n507) );
  BUFX3 aes_core_sbox_inst_U1563 ( .A(aes_core_sbox_inst_n507), .Y(
        aes_core_sbox_inst_n66) );
  NOR2X1 aes_core_sbox_inst_U1562 ( .A(aes_core_sbox_inst_n15), .B(
        aes_core_n29), .Y(aes_core_sbox_inst_n774) );
  BUFX3 aes_core_sbox_inst_U1561 ( .A(aes_core_sbox_inst_n774), .Y(
        aes_core_sbox_inst_n106) );
  NOR2X1 aes_core_sbox_inst_U1560 ( .A(aes_core_n5), .B(aes_core_n6), .Y(
        aes_core_sbox_inst_n479) );
  BUFX3 aes_core_sbox_inst_U1559 ( .A(aes_core_sbox_inst_n479), .Y(
        aes_core_sbox_inst_n71) );
  OAI221X1 aes_core_sbox_inst_U1558 ( .A0(aes_core_sbox_inst_n144), .A1(
        aes_core_sbox_inst_n1637), .B0(aes_core_sbox_inst_n57), .B1(
        aes_core_sbox_inst_n1654), .C0(aes_core_sbox_inst_n1640), .Y(
        aes_core_sbox_inst_n1396) );
  INVX1 aes_core_sbox_inst_U1557 ( .A(aes_core_sbox_inst_n342), .Y(
        aes_core_sbox_inst_n1647) );
  AOI211X1 aes_core_sbox_inst_U1556 ( .A0(aes_core_sbox_inst_n1395), .A1(
        aes_core_sbox_inst_n34), .B0(aes_core_sbox_inst_n1396), .C0(
        aes_core_sbox_inst_n1647), .Y(aes_core_sbox_inst_n1394) );
  OAI22X1 aes_core_sbox_inst_U1555 ( .A0(aes_core_sbox_inst_n1623), .A1(
        aes_core_sbox_inst_n370), .B0(aes_core_sbox_inst_n1394), .B1(
        aes_core_sbox_inst_n1621), .Y(aes_core_sbox_inst_n1389) );
  INVX1 aes_core_sbox_inst_U1554 ( .A(aes_core_sbox_inst_n476), .Y(
        aes_core_sbox_inst_n1710) );
  AOI211X1 aes_core_sbox_inst_U1553 ( .A0(aes_core_sbox_inst_n71), .A1(
        aes_core_sbox_inst_n1730), .B0(aes_core_sbox_inst_n480), .C0(
        aes_core_sbox_inst_n481), .Y(aes_core_sbox_inst_n473) );
  AOI211X1 aes_core_sbox_inst_U1552 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n1731), .B0(aes_core_sbox_inst_n475), .C0(
        aes_core_sbox_inst_n1710), .Y(aes_core_sbox_inst_n474) );
  OAI22X1 aes_core_sbox_inst_U1551 ( .A0(aes_core_sbox_inst_n56), .A1(
        aes_core_sbox_inst_n473), .B0(aes_core_sbox_inst_n474), .B1(
        aes_core_sbox_inst_n1684), .Y(aes_core_sbox_inst_n465) );
  INVX1 aes_core_sbox_inst_U1550 ( .A(aes_core_sbox_inst_n1071), .Y(
        aes_core_sbox_inst_n1592) );
  AOI211X1 aes_core_sbox_inst_U1549 ( .A0(aes_core_sbox_inst_n97), .A1(
        aes_core_sbox_inst_n1612), .B0(aes_core_sbox_inst_n1075), .C0(
        aes_core_sbox_inst_n1076), .Y(aes_core_sbox_inst_n1068) );
  AOI211X1 aes_core_sbox_inst_U1548 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n1613), .B0(aes_core_sbox_inst_n1070), .C0(
        aes_core_sbox_inst_n1592), .Y(aes_core_sbox_inst_n1069) );
  OAI22X1 aes_core_sbox_inst_U1547 ( .A0(aes_core_sbox_inst_n62), .A1(
        aes_core_sbox_inst_n1068), .B0(aes_core_sbox_inst_n1069), .B1(
        aes_core_sbox_inst_n1566), .Y(aes_core_sbox_inst_n1060) );
  INVX1 aes_core_sbox_inst_U1546 ( .A(aes_core_sbox_inst_n709), .Y(
        aes_core_sbox_inst_n233) );
  AOI211X1 aes_core_sbox_inst_U1545 ( .A0(aes_core_sbox_inst_n110), .A1(
        aes_core_sbox_inst_n253), .B0(aes_core_sbox_inst_n713), .C0(
        aes_core_sbox_inst_n714), .Y(aes_core_sbox_inst_n706) );
  AOI211X1 aes_core_sbox_inst_U1544 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n254), .B0(aes_core_sbox_inst_n708), .C0(
        aes_core_sbox_inst_n233), .Y(aes_core_sbox_inst_n707) );
  OAI22X1 aes_core_sbox_inst_U1543 ( .A0(aes_core_sbox_inst_n64), .A1(
        aes_core_sbox_inst_n706), .B0(aes_core_sbox_inst_n707), .B1(
        aes_core_sbox_inst_n208), .Y(aes_core_sbox_inst_n698) );
  AOI21X1 aes_core_sbox_inst_U1542 ( .A0(aes_core_sbox_inst_n1705), .A1(
        aes_core_sbox_inst_n518), .B0(aes_core_sbox_inst_n48), .Y(
        aes_core_sbox_inst_n525) );
  AOI21X1 aes_core_sbox_inst_U1541 ( .A0(aes_core_sbox_inst_n1587), .A1(
        aes_core_sbox_inst_n1113), .B0(aes_core_sbox_inst_n21), .Y(
        aes_core_sbox_inst_n1120) );
  AOI21X1 aes_core_sbox_inst_U1540 ( .A0(aes_core_sbox_inst_n228), .A1(
        aes_core_sbox_inst_n785), .B0(aes_core_sbox_inst_n13), .Y(
        aes_core_sbox_inst_n792) );
  AOI31X1 aes_core_sbox_inst_U1539 ( .A0(aes_core_n30), .A1(
        aes_core_sbox_inst_n259), .A2(aes_core_sbox_inst_n721), .B0(
        aes_core_sbox_inst_n792), .Y(aes_core_sbox_inst_n786) );
  AOI21X1 aes_core_sbox_inst_U1538 ( .A0(aes_core_sbox_inst_n58), .A1(
        aes_core_sbox_inst_n86), .B0(aes_core_sbox_inst_n1342), .Y(
        aes_core_sbox_inst_n1341) );
  AOI31X1 aes_core_sbox_inst_U1537 ( .A0(aes_core_sbox_inst_n1339), .A1(
        aes_core_sbox_inst_n1340), .A2(aes_core_sbox_inst_n1341), .B0(
        aes_core_sbox_inst_n182), .Y(aes_core_sbox_inst_n1338) );
  AOI2BB2X1 aes_core_sbox_inst_U1536 ( .B0(aes_core_sbox_inst_n401), .B1(
        aes_core_sbox_inst_n65), .A0N(aes_core_sbox_inst_n403), .A1N(
        aes_core_sbox_inst_n139), .Y(aes_core_sbox_inst_n388) );
  AOI221X1 aes_core_sbox_inst_U1535 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n192), .B0(aes_core_sbox_inst_n392), .B1(
        aes_core_sbox_inst_n128), .C0(aes_core_sbox_inst_n393), .Y(
        aes_core_sbox_inst_n390) );
  AOI31X1 aes_core_sbox_inst_U1534 ( .A0(aes_core_sbox_inst_n52), .A1(
        aes_core_sbox_inst_n50), .A2(aes_core_sbox_inst_n399), .B0(
        aes_core_sbox_inst_n400), .Y(aes_core_sbox_inst_n389) );
  AOI31X1 aes_core_sbox_inst_U1533 ( .A0(aes_core_sbox_inst_n388), .A1(
        aes_core_sbox_inst_n389), .A2(aes_core_sbox_inst_n390), .B0(
        aes_core_sbox_inst_n56), .Y(aes_core_sbox_inst_n376) );
  AOI2BB2X1 aes_core_sbox_inst_U1532 ( .B0(aes_core_sbox_inst_n996), .B1(
        aes_core_sbox_inst_n91), .A0N(aes_core_sbox_inst_n998), .A1N(
        aes_core_sbox_inst_n130), .Y(aes_core_sbox_inst_n983) );
  AOI221X1 aes_core_sbox_inst_U1531 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n170), .B0(aes_core_sbox_inst_n987), .B1(
        aes_core_sbox_inst_n123), .C0(aes_core_sbox_inst_n988), .Y(
        aes_core_sbox_inst_n985) );
  AOI31X1 aes_core_sbox_inst_U1530 ( .A0(aes_core_sbox_inst_n28), .A1(
        aes_core_sbox_inst_n25), .A2(aes_core_sbox_inst_n994), .B0(
        aes_core_sbox_inst_n995), .Y(aes_core_sbox_inst_n984) );
  AOI31X1 aes_core_sbox_inst_U1529 ( .A0(aes_core_sbox_inst_n983), .A1(
        aes_core_sbox_inst_n984), .A2(aes_core_sbox_inst_n985), .B0(
        aes_core_sbox_inst_n62), .Y(aes_core_sbox_inst_n971) );
  AOI2BB2X1 aes_core_sbox_inst_U1528 ( .B0(aes_core_sbox_inst_n634), .B1(
        aes_core_sbox_inst_n105), .A0N(aes_core_sbox_inst_n636), .A1N(
        aes_core_sbox_inst_n135), .Y(aes_core_sbox_inst_n621) );
  AOI221X1 aes_core_sbox_inst_U1527 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n154), .B0(aes_core_sbox_inst_n625), .B1(
        aes_core_sbox_inst_n119), .C0(aes_core_sbox_inst_n626), .Y(
        aes_core_sbox_inst_n623) );
  AOI31X1 aes_core_sbox_inst_U1526 ( .A0(aes_core_sbox_inst_n19), .A1(
        aes_core_sbox_inst_n17), .A2(aes_core_sbox_inst_n632), .B0(
        aes_core_sbox_inst_n633), .Y(aes_core_sbox_inst_n622) );
  AOI31X1 aes_core_sbox_inst_U1525 ( .A0(aes_core_sbox_inst_n621), .A1(
        aes_core_sbox_inst_n622), .A2(aes_core_sbox_inst_n623), .B0(
        aes_core_sbox_inst_n64), .Y(aes_core_sbox_inst_n609) );
  AOI221X1 aes_core_sbox_inst_U1524 ( .A0(aes_core_sbox_inst_n90), .A1(
        aes_core_sbox_inst_n58), .B0(aes_core_sbox_inst_n307), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n1338), .Y(
        aes_core_sbox_inst_n1337) );
  AOI2BB2X1 aes_core_sbox_inst_U1523 ( .B0(aes_core_sbox_inst_n1344), .B1(
        aes_core_sbox_inst_n87), .A0N(aes_core_sbox_inst_n1345), .A1N(
        aes_core_sbox_inst_n143), .Y(aes_core_sbox_inst_n1335) );
  AOI31X1 aes_core_sbox_inst_U1522 ( .A0(aes_core_sbox_inst_n81), .A1(
        aes_core_sbox_inst_n38), .A2(aes_core_sbox_inst_n359), .B0(
        aes_core_sbox_inst_n1343), .Y(aes_core_sbox_inst_n1336) );
  AOI31X1 aes_core_sbox_inst_U1521 ( .A0(aes_core_sbox_inst_n1335), .A1(
        aes_core_sbox_inst_n1336), .A2(aes_core_sbox_inst_n1337), .B0(
        aes_core_n16), .Y(aes_core_sbox_inst_n1328) );
  AOI31X1 aes_core_sbox_inst_U1520 ( .A0(aes_core_sbox_inst_n57), .A1(
        aes_core_n14), .A2(aes_core_sbox_inst_n359), .B0(
        aes_core_sbox_inst_n1627), .Y(aes_core_sbox_inst_n1475) );
  NAND3X1 aes_core_sbox_inst_U1519 ( .A(aes_core_sbox_inst_n58), .B(
        aes_core_sbox_inst_n1656), .C(aes_core_sbox_inst_n293), .Y(
        aes_core_sbox_inst_n1476) );
  AOI22X1 aes_core_sbox_inst_U1518 ( .A0(aes_core_sbox_inst_n57), .A1(
        aes_core_sbox_inst_n1333), .B0(aes_core_sbox_inst_n89), .B1(
        aes_core_sbox_inst_n80), .Y(aes_core_sbox_inst_n1332) );
  AOI31X1 aes_core_sbox_inst_U1517 ( .A0(aes_core_sbox_inst_n59), .A1(
        aes_core_sbox_inst_n33), .A2(aes_core_sbox_inst_n143), .B0(
        aes_core_sbox_inst_n277), .Y(aes_core_sbox_inst_n1330) );
  NAND3BX1 aes_core_sbox_inst_U1516 ( .AN(aes_core_sbox_inst_n1334), .B(
        aes_core_sbox_inst_n124), .C(aes_core_n14), .Y(
        aes_core_sbox_inst_n1331) );
  AOI31X1 aes_core_sbox_inst_U1515 ( .A0(aes_core_sbox_inst_n1330), .A1(
        aes_core_sbox_inst_n1331), .A2(aes_core_sbox_inst_n1332), .B0(
        aes_core_sbox_inst_n1622), .Y(aes_core_sbox_inst_n1329) );
  AOI31X1 aes_core_sbox_inst_U1514 ( .A0(aes_core_n6), .A1(
        aes_core_sbox_inst_n1727), .A2(aes_core_sbox_inst_n70), .B0(
        aes_core_sbox_inst_n387), .Y(aes_core_sbox_inst_n378) );
  AOI22X1 aes_core_sbox_inst_U1513 ( .A0(aes_core_sbox_inst_n199), .A1(
        aes_core_sbox_inst_n381), .B0(aes_core_sbox_inst_n76), .B1(
        aes_core_sbox_inst_n6), .Y(aes_core_sbox_inst_n380) );
  NAND3X1 aes_core_sbox_inst_U1512 ( .A(aes_core_sbox_inst_n138), .B(
        aes_core_sbox_inst_n55), .C(aes_core_sbox_inst_n385), .Y(
        aes_core_sbox_inst_n379) );
  AOI31X1 aes_core_sbox_inst_U1511 ( .A0(aes_core_sbox_inst_n378), .A1(
        aes_core_sbox_inst_n379), .A2(aes_core_sbox_inst_n380), .B0(
        aes_core_sbox_inst_n1684), .Y(aes_core_sbox_inst_n377) );
  AOI31X1 aes_core_sbox_inst_U1510 ( .A0(aes_core_sbox_inst_n61), .A1(
        aes_core_sbox_inst_n1609), .A2(aes_core_sbox_inst_n96), .B0(
        aes_core_sbox_inst_n982), .Y(aes_core_sbox_inst_n973) );
  AOI22X1 aes_core_sbox_inst_U1509 ( .A0(aes_core_sbox_inst_n174), .A1(
        aes_core_sbox_inst_n976), .B0(aes_core_sbox_inst_n102), .B1(
        aes_core_sbox_inst_n7), .Y(aes_core_sbox_inst_n975) );
  NAND3X1 aes_core_sbox_inst_U1508 ( .A(aes_core_sbox_inst_n129), .B(
        aes_core_sbox_inst_n60), .C(aes_core_sbox_inst_n980), .Y(
        aes_core_sbox_inst_n974) );
  AOI31X1 aes_core_sbox_inst_U1507 ( .A0(aes_core_sbox_inst_n973), .A1(
        aes_core_sbox_inst_n974), .A2(aes_core_sbox_inst_n975), .B0(
        aes_core_sbox_inst_n1566), .Y(aes_core_sbox_inst_n972) );
  AOI31X1 aes_core_sbox_inst_U1506 ( .A0(aes_core_n30), .A1(
        aes_core_sbox_inst_n250), .A2(aes_core_sbox_inst_n109), .B0(
        aes_core_sbox_inst_n620), .Y(aes_core_sbox_inst_n611) );
  AOI22X1 aes_core_sbox_inst_U1505 ( .A0(aes_core_sbox_inst_n159), .A1(
        aes_core_sbox_inst_n614), .B0(aes_core_sbox_inst_n114), .B1(
        aes_core_sbox_inst_n616), .Y(aes_core_sbox_inst_n613) );
  NAND3X1 aes_core_sbox_inst_U1504 ( .A(aes_core_sbox_inst_n134), .B(
        aes_core_sbox_inst_n63), .C(aes_core_sbox_inst_n618), .Y(
        aes_core_sbox_inst_n612) );
  AOI31X1 aes_core_sbox_inst_U1503 ( .A0(aes_core_sbox_inst_n611), .A1(
        aes_core_sbox_inst_n612), .A2(aes_core_sbox_inst_n613), .B0(
        aes_core_sbox_inst_n208), .Y(aes_core_sbox_inst_n610) );
  OAI32X1 aes_core_sbox_inst_U1502 ( .A0(aes_core_sbox_inst_n1704), .A1(
        aes_core_sbox_inst_n55), .A2(aes_core_sbox_inst_n53), .B0(
        aes_core_sbox_inst_n126), .B1(aes_core_sbox_inst_n1700), .Y(
        aes_core_sbox_inst_n533) );
  AOI21X1 aes_core_sbox_inst_U1501 ( .A0(aes_core_sbox_inst_n78), .A1(
        aes_core_sbox_inst_n6), .B0(aes_core_sbox_inst_n533), .Y(
        aes_core_sbox_inst_n532) );
  OAI211X1 aes_core_sbox_inst_U1500 ( .A0(aes_core_sbox_inst_n1718), .A1(
        aes_core_sbox_inst_n141), .B0(aes_core_sbox_inst_n459), .C0(
        aes_core_sbox_inst_n532), .Y(aes_core_sbox_inst_n531) );
  OAI32X1 aes_core_sbox_inst_U1499 ( .A0(aes_core_sbox_inst_n1586), .A1(
        aes_core_sbox_inst_n60), .A2(aes_core_sbox_inst_n29), .B0(
        aes_core_sbox_inst_n121), .B1(aes_core_sbox_inst_n1582), .Y(
        aes_core_sbox_inst_n1128) );
  AOI21X1 aes_core_sbox_inst_U1498 ( .A0(aes_core_sbox_inst_n104), .A1(
        aes_core_sbox_inst_n7), .B0(aes_core_sbox_inst_n1128), .Y(
        aes_core_sbox_inst_n1127) );
  OAI211X1 aes_core_sbox_inst_U1497 ( .A0(aes_core_sbox_inst_n1600), .A1(
        aes_core_sbox_inst_n132), .B0(aes_core_sbox_inst_n1054), .C0(
        aes_core_sbox_inst_n1127), .Y(aes_core_sbox_inst_n1126) );
  OAI32X1 aes_core_sbox_inst_U1496 ( .A0(aes_core_sbox_inst_n227), .A1(
        aes_core_sbox_inst_n63), .A2(aes_core_sbox_inst_n19), .B0(
        aes_core_sbox_inst_n117), .B1(aes_core_sbox_inst_n11), .Y(
        aes_core_sbox_inst_n800) );
  AOI21X1 aes_core_sbox_inst_U1495 ( .A0(aes_core_sbox_inst_n116), .A1(
        aes_core_sbox_inst_n8), .B0(aes_core_sbox_inst_n800), .Y(
        aes_core_sbox_inst_n799) );
  OAI211X1 aes_core_sbox_inst_U1494 ( .A0(aes_core_sbox_inst_n16), .A1(
        aes_core_sbox_inst_n1), .B0(aes_core_sbox_inst_n692), .C0(
        aes_core_sbox_inst_n799), .Y(aes_core_sbox_inst_n798) );
  OAI211X1 aes_core_sbox_inst_U1493 ( .A0(aes_core_sbox_inst_n162), .A1(
        aes_core_sbox_inst_n219), .B0(aes_core_sbox_inst_n959), .C0(
        aes_core_sbox_inst_n960), .Y(aes_core_sbox_inst_n952) );
  OAI222X1 aes_core_sbox_inst_U1492 ( .A0(aes_core_sbox_inst_n937), .A1(
        aes_core_sbox_inst_n209), .B0(aes_core_sbox_inst_n938), .B1(
        aes_core_sbox_inst_n208), .C0(aes_core_sbox_inst_n64), .C1(
        aes_core_sbox_inst_n939), .Y(aes_core_sbox_inst_n936) );
  AOI22X1 aes_core_sbox_inst_U1491 ( .A0(aes_core_sbox_inst_n64), .A1(
        aes_core_sbox_inst_n952), .B0(aes_core_sbox_inst_n953), .B1(
        aes_core_sbox_inst_n209), .Y(aes_core_sbox_inst_n935) );
  OAI2BB2X1 aes_core_sbox_inst_U1490 ( .B0(aes_core_n33), .B1(
        aes_core_sbox_inst_n935), .A0N(aes_core_n33), .A1N(
        aes_core_sbox_inst_n936), .Y(aes_core_new_sboxw[24]) );
  AOI221X1 aes_core_sbox_inst_U1489 ( .A0(aes_core_sbox_inst_n78), .A1(
        aes_core_sbox_inst_n54), .B0(aes_core_sbox_inst_n77), .B1(
        aes_core_sbox_inst_n197), .C0(aes_core_sbox_inst_n1551), .Y(
        aes_core_sbox_inst_n1550) );
  NAND4BX1 aes_core_sbox_inst_U1488 ( .AN(aes_core_sbox_inst_n421), .B(
        aes_core_sbox_inst_n1706), .C(aes_core_sbox_inst_n1549), .D(
        aes_core_sbox_inst_n1550), .Y(aes_core_sbox_inst_n1546) );
  NOR3X1 aes_core_sbox_inst_U1487 ( .A(aes_core_sbox_inst_n126), .B(
        aes_core_n5), .C(aes_core_sbox_inst_n48), .Y(aes_core_sbox_inst_n1548)
         );
  AOI211X1 aes_core_sbox_inst_U1486 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n1546), .B0(aes_core_sbox_inst_n1547), .C0(
        aes_core_sbox_inst_n1548), .Y(aes_core_sbox_inst_n1537) );
  AOI221X1 aes_core_sbox_inst_U1485 ( .A0(aes_core_sbox_inst_n104), .A1(
        aes_core_sbox_inst_n30), .B0(aes_core_sbox_inst_n103), .B1(
        aes_core_sbox_inst_n174), .C0(aes_core_sbox_inst_n1309), .Y(
        aes_core_sbox_inst_n1308) );
  NAND4BX1 aes_core_sbox_inst_U1484 ( .AN(aes_core_sbox_inst_n1016), .B(
        aes_core_sbox_inst_n1588), .C(aes_core_sbox_inst_n1307), .D(
        aes_core_sbox_inst_n1308), .Y(aes_core_sbox_inst_n1304) );
  NOR3X1 aes_core_sbox_inst_U1483 ( .A(aes_core_sbox_inst_n121), .B(
        aes_core_n21), .C(aes_core_sbox_inst_n21), .Y(aes_core_sbox_inst_n1306) );
  AOI211X1 aes_core_sbox_inst_U1482 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1304), .B0(aes_core_sbox_inst_n1305), .C0(
        aes_core_sbox_inst_n1306), .Y(aes_core_sbox_inst_n1295) );
  AOI221X1 aes_core_sbox_inst_U1481 ( .A0(aes_core_sbox_inst_n116), .A1(
        aes_core_sbox_inst_n259), .B0(aes_core_sbox_inst_n115), .B1(
        aes_core_sbox_inst_n160), .C0(aes_core_sbox_inst_n951), .Y(
        aes_core_sbox_inst_n950) );
  NAND4BX1 aes_core_sbox_inst_U1480 ( .AN(aes_core_sbox_inst_n654), .B(
        aes_core_sbox_inst_n229), .C(aes_core_sbox_inst_n949), .D(
        aes_core_sbox_inst_n950), .Y(aes_core_sbox_inst_n946) );
  NOR3X1 aes_core_sbox_inst_U1479 ( .A(aes_core_sbox_inst_n117), .B(
        aes_core_n29), .C(aes_core_sbox_inst_n13), .Y(aes_core_sbox_inst_n948)
         );
  AOI211X1 aes_core_sbox_inst_U1478 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n946), .B0(aes_core_sbox_inst_n947), .C0(
        aes_core_sbox_inst_n948), .Y(aes_core_sbox_inst_n937) );
  AOI31X1 aes_core_sbox_inst_U1477 ( .A0(aes_core_sbox_inst_n142), .A1(
        aes_core_n14), .A2(aes_core_sbox_inst_n359), .B0(
        aes_core_sbox_inst_n1634), .Y(aes_core_sbox_inst_n361) );
  AOI221X1 aes_core_sbox_inst_U1476 ( .A0(aes_core_sbox_inst_n1379), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n1380), .B1(
        aes_core_sbox_inst_n47), .C0(aes_core_sbox_inst_n346), .Y(
        aes_core_sbox_inst_n1378) );
  OAI221X1 aes_core_sbox_inst_U1475 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n1654), .B0(aes_core_sbox_inst_n58), .B1(
        aes_core_sbox_inst_n1638), .C0(aes_core_sbox_inst_n1378), .Y(
        aes_core_sbox_inst_n1373) );
  OAI211X1 aes_core_sbox_inst_U1474 ( .A0(aes_core_sbox_inst_n58), .A1(
        aes_core_sbox_inst_n1651), .B0(aes_core_sbox_inst_n1640), .C0(
        aes_core_sbox_inst_n1514), .Y(aes_core_sbox_inst_n1510) );
  AND3X2 aes_core_sbox_inst_U1473 ( .A(aes_core_sbox_inst_n625), .B(
        aes_core_sbox_inst_n1), .C(aes_core_sbox_inst_n64), .Y(
        aes_core_sbox_inst_n920) );
  AOI222X1 aes_core_sbox_inst_U1472 ( .A0(aes_core_sbox_inst_n907), .A1(
        aes_core_sbox_inst_n209), .B0(aes_core_sbox_inst_n607), .B1(
        aes_core_sbox_inst_n908), .C0(aes_core_sbox_inst_n859), .C1(
        aes_core_sbox_inst_n909), .Y(aes_core_sbox_inst_n906) );
  NOR4BX1 aes_core_sbox_inst_U1471 ( .AN(aes_core_sbox_inst_n919), .B(
        aes_core_sbox_inst_n920), .C(aes_core_sbox_inst_n921), .D(
        aes_core_sbox_inst_n922), .Y(aes_core_sbox_inst_n905) );
  OAI22X1 aes_core_sbox_inst_U1470 ( .A0(aes_core_sbox_inst_n905), .A1(
        aes_core_sbox_inst_n206), .B0(aes_core_n33), .B1(
        aes_core_sbox_inst_n906), .Y(aes_core_new_sboxw[25]) );
  AOI21X1 aes_core_sbox_inst_U1469 ( .A0(aes_core_sbox_inst_n1241), .A1(
        aes_core_sbox_inst_n1242), .B0(aes_core_n25), .Y(
        aes_core_sbox_inst_n1231) );
  NAND4X1 aes_core_sbox_inst_U1468 ( .A(aes_core_sbox_inst_n1256), .B(
        aes_core_sbox_inst_n1257), .C(aes_core_sbox_inst_n1258), .D(
        aes_core_sbox_inst_n1259), .Y(aes_core_sbox_inst_n1230) );
  AOI211X1 aes_core_sbox_inst_U1467 ( .A0(aes_core_sbox_inst_n1197), .A1(
        aes_core_sbox_inst_n1230), .B0(aes_core_sbox_inst_n1231), .C0(
        aes_core_sbox_inst_n1232), .Y(aes_core_sbox_inst_n1229) );
  INVX1 aes_core_sbox_inst_U1466 ( .A(aes_core_sbox_inst_n1229), .Y(
        aes_core_new_sboxw[18]) );
  AOI21X1 aes_core_sbox_inst_U1465 ( .A0(aes_core_sbox_inst_n1515), .A1(
        aes_core_sbox_inst_n1516), .B0(aes_core_n17), .Y(
        aes_core_sbox_inst_n1506) );
  NAND4X1 aes_core_sbox_inst_U1464 ( .A(aes_core_sbox_inst_n1429), .B(
        aes_core_sbox_inst_n360), .C(aes_core_sbox_inst_n1530), .D(
        aes_core_sbox_inst_n1531), .Y(aes_core_sbox_inst_n1505) );
  AOI211X1 aes_core_sbox_inst_U1463 ( .A0(aes_core_sbox_inst_n1478), .A1(
        aes_core_sbox_inst_n1505), .B0(aes_core_sbox_inst_n1506), .C0(
        aes_core_sbox_inst_n1507), .Y(aes_core_sbox_inst_n1504) );
  INVX1 aes_core_sbox_inst_U1462 ( .A(aes_core_sbox_inst_n1504), .Y(
        aes_core_new_sboxw[10]) );
  AOI21X1 aes_core_sbox_inst_U1461 ( .A0(aes_core_sbox_inst_n736), .A1(
        aes_core_sbox_inst_n737), .B0(aes_core_n9), .Y(aes_core_sbox_inst_n726) );
  NAND4X1 aes_core_sbox_inst_U1460 ( .A(aes_core_sbox_inst_n751), .B(
        aes_core_sbox_inst_n752), .C(aes_core_sbox_inst_n753), .D(
        aes_core_sbox_inst_n754), .Y(aes_core_sbox_inst_n725) );
  AOI211X1 aes_core_sbox_inst_U1459 ( .A0(aes_core_sbox_inst_n572), .A1(
        aes_core_sbox_inst_n725), .B0(aes_core_sbox_inst_n726), .C0(
        aes_core_sbox_inst_n727), .Y(aes_core_sbox_inst_n724) );
  INVX1 aes_core_sbox_inst_U1458 ( .A(aes_core_sbox_inst_n724), .Y(
        aes_core_new_sboxw[2]) );
  NAND4BX1 aes_core_sbox_inst_U1457 ( .AN(aes_core_sbox_inst_n1423), .B(
        aes_core_sbox_inst_n1484), .C(aes_core_sbox_inst_n1499), .D(
        aes_core_sbox_inst_n1500), .Y(aes_core_sbox_inst_n1472) );
  AOI21X1 aes_core_sbox_inst_U1456 ( .A0(aes_core_sbox_inst_n1485), .A1(
        aes_core_sbox_inst_n1486), .B0(aes_core_n17), .Y(
        aes_core_sbox_inst_n1473) );
  AOI211X1 aes_core_sbox_inst_U1455 ( .A0(aes_core_sbox_inst_n1471), .A1(
        aes_core_sbox_inst_n1472), .B0(aes_core_sbox_inst_n1473), .C0(
        aes_core_sbox_inst_n1474), .Y(aes_core_sbox_inst_n1470) );
  INVX1 aes_core_sbox_inst_U1454 ( .A(aes_core_sbox_inst_n1470), .Y(
        aes_core_new_sboxw[11]) );
  AOI21X1 aes_core_sbox_inst_U1453 ( .A0(aes_core_sbox_inst_n677), .A1(
        aes_core_sbox_inst_n678), .B0(aes_core_sbox_inst_n211), .Y(
        aes_core_sbox_inst_n676) );
  AOI211X1 aes_core_sbox_inst_U1452 ( .A0(aes_core_sbox_inst_n697), .A1(
        aes_core_sbox_inst_n64), .B0(aes_core_sbox_inst_n698), .C0(
        aes_core_sbox_inst_n699), .Y(aes_core_sbox_inst_n671) );
  AOI211X1 aes_core_sbox_inst_U1451 ( .A0(aes_core_sbox_inst_n673), .A1(
        aes_core_sbox_inst_n674), .B0(aes_core_sbox_inst_n675), .C0(
        aes_core_sbox_inst_n676), .Y(aes_core_sbox_inst_n672) );
  OAI22X1 aes_core_sbox_inst_U1450 ( .A0(aes_core_n33), .A1(
        aes_core_sbox_inst_n671), .B0(aes_core_sbox_inst_n672), .B1(
        aes_core_sbox_inst_n206), .Y(aes_core_new_sboxw[30]) );
  AOI211X1 aes_core_sbox_inst_U1449 ( .A0(aes_core_sbox_inst_n90), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n1430), .C0(
        aes_core_sbox_inst_n1431), .Y(aes_core_sbox_inst_n1427) );
  AOI32X1 aes_core_sbox_inst_U1448 ( .A0(aes_core_sbox_inst_n1656), .A1(
        aes_core_sbox_inst_n144), .A2(aes_core_sbox_inst_n359), .B0(
        aes_core_sbox_inst_n1631), .B1(aes_core_sbox_inst_n57), .Y(
        aes_core_sbox_inst_n1428) );
  AOI222X1 aes_core_sbox_inst_U1447 ( .A0(aes_core_sbox_inst_n87), .A1(
        aes_core_sbox_inst_n44), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n321), .C0(aes_core_sbox_inst_n79), .C1(
        aes_core_sbox_inst_n85), .Y(aes_core_sbox_inst_n1426) );
  OAI221X1 aes_core_sbox_inst_U1446 ( .A0(aes_core_sbox_inst_n1426), .A1(
        aes_core_sbox_inst_n31), .B0(aes_core_sbox_inst_n1427), .B1(
        aes_core_sbox_inst_n181), .C0(aes_core_sbox_inst_n1428), .Y(
        aes_core_sbox_inst_n1415) );
  AOI211X1 aes_core_sbox_inst_U1445 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n43), .B0(aes_core_sbox_inst_n1453), .C0(
        aes_core_sbox_inst_n1454), .Y(aes_core_sbox_inst_n1452) );
  AOI211X1 aes_core_sbox_inst_U1444 ( .A0(aes_core_sbox_inst_n367), .A1(
        aes_core_sbox_inst_n57), .B0(aes_core_sbox_inst_n1456), .C0(
        aes_core_sbox_inst_n356), .Y(aes_core_sbox_inst_n1450) );
  AOI21X1 aes_core_sbox_inst_U1443 ( .A0(aes_core_sbox_inst_n85), .A1(
        aes_core_sbox_inst_n1678), .B0(aes_core_sbox_inst_n1363), .Y(
        aes_core_sbox_inst_n1451) );
  OAI222X1 aes_core_sbox_inst_U1442 ( .A0(aes_core_sbox_inst_n1450), .A1(
        aes_core_sbox_inst_n181), .B0(aes_core_sbox_inst_n1451), .B1(
        aes_core_sbox_inst_n1630), .C0(aes_core_sbox_inst_n184), .C1(
        aes_core_sbox_inst_n1452), .Y(aes_core_sbox_inst_n1441) );
  AOI221X1 aes_core_sbox_inst_U1441 ( .A0(aes_core_sbox_inst_n10), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n1333), .B1(
        aes_core_sbox_inst_n44), .C0(aes_core_sbox_inst_n1425), .Y(
        aes_core_sbox_inst_n1503) );
  AOI22X1 aes_core_sbox_inst_U1440 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n90), .B1(
        aes_core_sbox_inst_n1678), .Y(aes_core_sbox_inst_n1502) );
  OAI211X1 aes_core_sbox_inst_U1439 ( .A0(aes_core_sbox_inst_n41), .A1(
        aes_core_sbox_inst_n32), .B0(aes_core_sbox_inst_n1502), .C0(
        aes_core_sbox_inst_n1503), .Y(aes_core_sbox_inst_n1501) );
  AOI222X1 aes_core_sbox_inst_U1438 ( .A0(aes_core_sbox_inst_n184), .A1(
        aes_core_sbox_inst_n1501), .B0(aes_core_sbox_inst_n1344), .B1(
        aes_core_sbox_inst_n82), .C0(aes_core_sbox_inst_n292), .C1(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n1500) );
  OAI211X1 aes_core_sbox_inst_U1437 ( .A0(aes_core_sbox_inst_n200), .A1(
        aes_core_sbox_inst_n1695), .B0(aes_core_sbox_inst_n1559), .C0(
        aes_core_sbox_inst_n1560), .Y(aes_core_sbox_inst_n1552) );
  OAI222X1 aes_core_sbox_inst_U1436 ( .A0(aes_core_sbox_inst_n1537), .A1(
        aes_core_sbox_inst_n1685), .B0(aes_core_sbox_inst_n1538), .B1(
        aes_core_sbox_inst_n1684), .C0(aes_core_sbox_inst_n56), .C1(
        aes_core_sbox_inst_n1539), .Y(aes_core_sbox_inst_n1536) );
  AOI22X1 aes_core_sbox_inst_U1435 ( .A0(aes_core_sbox_inst_n56), .A1(
        aes_core_sbox_inst_n1552), .B0(aes_core_sbox_inst_n1553), .B1(
        aes_core_sbox_inst_n1685), .Y(aes_core_sbox_inst_n1535) );
  OAI2BB2X1 aes_core_sbox_inst_U1434 ( .B0(aes_core_n9), .B1(
        aes_core_sbox_inst_n1535), .A0N(aes_core_n9), .A1N(
        aes_core_sbox_inst_n1536), .Y(aes_core_new_sboxw[0]) );
  OAI211X1 aes_core_sbox_inst_U1433 ( .A0(aes_core_sbox_inst_n175), .A1(
        aes_core_sbox_inst_n1577), .B0(aes_core_sbox_inst_n1317), .C0(
        aes_core_sbox_inst_n1318), .Y(aes_core_sbox_inst_n1310) );
  OAI222X1 aes_core_sbox_inst_U1432 ( .A0(aes_core_sbox_inst_n1295), .A1(
        aes_core_sbox_inst_n1567), .B0(aes_core_sbox_inst_n1296), .B1(
        aes_core_sbox_inst_n1566), .C0(aes_core_sbox_inst_n62), .C1(
        aes_core_sbox_inst_n1297), .Y(aes_core_sbox_inst_n1294) );
  AOI22X1 aes_core_sbox_inst_U1431 ( .A0(aes_core_sbox_inst_n62), .A1(
        aes_core_sbox_inst_n1310), .B0(aes_core_sbox_inst_n1311), .B1(
        aes_core_sbox_inst_n1567), .Y(aes_core_sbox_inst_n1293) );
  OAI2BB2X1 aes_core_sbox_inst_U1430 ( .B0(aes_core_n25), .B1(
        aes_core_sbox_inst_n1293), .A0N(aes_core_n25), .A1N(
        aes_core_sbox_inst_n1294), .Y(aes_core_new_sboxw[16]) );
  AOI22X1 aes_core_sbox_inst_U1429 ( .A0(aes_core_n16), .A1(
        aes_core_sbox_inst_n347), .B0(aes_core_sbox_inst_n348), .B1(
        aes_core_sbox_inst_n1623), .Y(aes_core_sbox_inst_n323) );
  NOR2X1 aes_core_sbox_inst_U1428 ( .A(aes_core_sbox_inst_n38), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n276) );
  AND3X2 aes_core_sbox_inst_U1427 ( .A(aes_core_sbox_inst_n987), .B(
        aes_core_sbox_inst_n133), .C(aes_core_sbox_inst_n62), .Y(
        aes_core_sbox_inst_n1278) );
  AOI222X1 aes_core_sbox_inst_U1426 ( .A0(aes_core_sbox_inst_n1265), .A1(
        aes_core_sbox_inst_n1567), .B0(aes_core_sbox_inst_n969), .B1(
        aes_core_sbox_inst_n1266), .C0(aes_core_sbox_inst_n1217), .C1(
        aes_core_sbox_inst_n1267), .Y(aes_core_sbox_inst_n1264) );
  NOR4BX1 aes_core_sbox_inst_U1425 ( .AN(aes_core_sbox_inst_n1277), .B(
        aes_core_sbox_inst_n1278), .C(aes_core_sbox_inst_n1279), .D(
        aes_core_sbox_inst_n1280), .Y(aes_core_sbox_inst_n1263) );
  OAI22X1 aes_core_sbox_inst_U1424 ( .A0(aes_core_sbox_inst_n1263), .A1(
        aes_core_sbox_inst_n450), .B0(aes_core_n25), .B1(
        aes_core_sbox_inst_n1264), .Y(aes_core_new_sboxw[17]) );
  AOI21X1 aes_core_sbox_inst_U1423 ( .A0(aes_core_sbox_inst_n1039), .A1(
        aes_core_sbox_inst_n1040), .B0(aes_core_sbox_inst_n1569), .Y(
        aes_core_sbox_inst_n1038) );
  AOI211X1 aes_core_sbox_inst_U1422 ( .A0(aes_core_sbox_inst_n1059), .A1(
        aes_core_sbox_inst_n62), .B0(aes_core_sbox_inst_n1060), .C0(
        aes_core_sbox_inst_n1061), .Y(aes_core_sbox_inst_n1033) );
  AOI211X1 aes_core_sbox_inst_U1421 ( .A0(aes_core_sbox_inst_n1035), .A1(
        aes_core_sbox_inst_n1036), .B0(aes_core_sbox_inst_n1037), .C0(
        aes_core_sbox_inst_n1038), .Y(aes_core_sbox_inst_n1034) );
  OAI22X1 aes_core_sbox_inst_U1420 ( .A0(aes_core_n25), .A1(
        aes_core_sbox_inst_n1033), .B0(aes_core_sbox_inst_n1034), .B1(
        aes_core_sbox_inst_n450), .Y(aes_core_new_sboxw[22]) );
  AND3X2 aes_core_sbox_inst_U1419 ( .A(aes_core_sbox_inst_n392), .B(
        aes_core_sbox_inst_n140), .C(aes_core_sbox_inst_n56), .Y(
        aes_core_sbox_inst_n1174) );
  AOI222X1 aes_core_sbox_inst_U1418 ( .A0(aes_core_sbox_inst_n1161), .A1(
        aes_core_sbox_inst_n1685), .B0(aes_core_sbox_inst_n374), .B1(
        aes_core_sbox_inst_n1162), .C0(aes_core_sbox_inst_n592), .C1(
        aes_core_sbox_inst_n1163), .Y(aes_core_sbox_inst_n1160) );
  NOR4BX1 aes_core_sbox_inst_U1417 ( .AN(aes_core_sbox_inst_n1173), .B(
        aes_core_sbox_inst_n1174), .C(aes_core_sbox_inst_n1175), .D(
        aes_core_sbox_inst_n1176), .Y(aes_core_sbox_inst_n1159) );
  OAI22X1 aes_core_sbox_inst_U1416 ( .A0(aes_core_sbox_inst_n1159), .A1(
        aes_core_sbox_inst_n1682), .B0(aes_core_n9), .B1(
        aes_core_sbox_inst_n1160), .Y(aes_core_new_sboxw[1]) );
  NAND4X1 aes_core_sbox_inst_U1415 ( .A(aes_core_sbox_inst_n1348), .B(
        aes_core_sbox_inst_n1638), .C(aes_core_sbox_inst_n1376), .D(
        aes_core_sbox_inst_n1377), .Y(aes_core_sbox_inst_n1375) );
  AOI211X1 aes_core_sbox_inst_U1414 ( .A0(aes_core_sbox_inst_n1388), .A1(
        aes_core_sbox_inst_n1623), .B0(aes_core_sbox_inst_n1389), .C0(
        aes_core_sbox_inst_n1390), .Y(aes_core_sbox_inst_n1369) );
  AOI222X1 aes_core_sbox_inst_U1413 ( .A0(aes_core_n16), .A1(
        aes_core_sbox_inst_n1371), .B0(aes_core_sbox_inst_n1372), .B1(
        aes_core_sbox_inst_n1373), .C0(aes_core_sbox_inst_n1374), .C1(
        aes_core_sbox_inst_n1375), .Y(aes_core_sbox_inst_n1370) );
  OAI22X1 aes_core_sbox_inst_U1412 ( .A0(aes_core_n17), .A1(
        aes_core_sbox_inst_n1369), .B0(aes_core_sbox_inst_n1370), .B1(
        aes_core_sbox_inst_n1620), .Y(aes_core_new_sboxw[14]) );
  AOI21X1 aes_core_sbox_inst_U1411 ( .A0(aes_core_sbox_inst_n444), .A1(
        aes_core_sbox_inst_n445), .B0(aes_core_sbox_inst_n1687), .Y(
        aes_core_sbox_inst_n443) );
  AOI211X1 aes_core_sbox_inst_U1410 ( .A0(aes_core_sbox_inst_n464), .A1(
        aes_core_sbox_inst_n56), .B0(aes_core_sbox_inst_n465), .C0(
        aes_core_sbox_inst_n466), .Y(aes_core_sbox_inst_n438) );
  AOI211X1 aes_core_sbox_inst_U1409 ( .A0(aes_core_sbox_inst_n440), .A1(
        aes_core_sbox_inst_n441), .B0(aes_core_sbox_inst_n442), .C0(
        aes_core_sbox_inst_n443), .Y(aes_core_sbox_inst_n439) );
  OAI22X1 aes_core_sbox_inst_U1408 ( .A0(aes_core_n9), .A1(
        aes_core_sbox_inst_n438), .B0(aes_core_sbox_inst_n439), .B1(
        aes_core_sbox_inst_n1682), .Y(aes_core_new_sboxw[6]) );
  AOI22X1 aes_core_sbox_inst_U1407 ( .A0(aes_core_sbox_inst_n64), .A1(
        aes_core_sbox_inst_n767), .B0(aes_core_sbox_inst_n768), .B1(
        aes_core_sbox_inst_n209), .Y(aes_core_sbox_inst_n759) );
  NOR4BBX1 aes_core_sbox_inst_U1406 ( .AN(aes_core_sbox_inst_n786), .BN(
        aes_core_sbox_inst_n787), .C(aes_core_sbox_inst_n633), .D(
        aes_core_sbox_inst_n620), .Y(aes_core_sbox_inst_n758) );
  AOI222X1 aes_core_sbox_inst_U1405 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n761), .B0(aes_core_sbox_inst_n762), .B1(
        aes_core_sbox_inst_n148), .C0(aes_core_sbox_inst_n637), .C1(
        aes_core_sbox_inst_n763), .Y(aes_core_sbox_inst_n760) );
  OAI222X1 aes_core_sbox_inst_U1404 ( .A0(aes_core_sbox_inst_n758), .A1(
        aes_core_sbox_inst_n205), .B0(aes_core_n33), .B1(
        aes_core_sbox_inst_n759), .C0(aes_core_sbox_inst_n760), .C1(
        aes_core_sbox_inst_n204), .Y(aes_core_new_sboxw[29]) );
  AOI22X1 aes_core_sbox_inst_U1403 ( .A0(aes_core_sbox_inst_n62), .A1(
        aes_core_sbox_inst_n1095), .B0(aes_core_sbox_inst_n1096), .B1(
        aes_core_sbox_inst_n1567), .Y(aes_core_sbox_inst_n1087) );
  NOR4BBX1 aes_core_sbox_inst_U1402 ( .AN(aes_core_sbox_inst_n1114), .BN(
        aes_core_sbox_inst_n1115), .C(aes_core_sbox_inst_n995), .D(
        aes_core_sbox_inst_n982), .Y(aes_core_sbox_inst_n1086) );
  AOI222X1 aes_core_sbox_inst_U1401 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1089), .B0(aes_core_sbox_inst_n1090), .B1(
        aes_core_sbox_inst_n167), .C0(aes_core_sbox_inst_n999), .C1(
        aes_core_sbox_inst_n1091), .Y(aes_core_sbox_inst_n1088) );
  OAI222X1 aes_core_sbox_inst_U1400 ( .A0(aes_core_sbox_inst_n1086), .A1(
        aes_core_sbox_inst_n316), .B0(aes_core_n25), .B1(
        aes_core_sbox_inst_n1087), .C0(aes_core_sbox_inst_n1088), .C1(
        aes_core_sbox_inst_n273), .Y(aes_core_new_sboxw[21]) );
  AOI22X1 aes_core_sbox_inst_U1399 ( .A0(aes_core_n16), .A1(
        aes_core_sbox_inst_n1415), .B0(aes_core_sbox_inst_n1416), .B1(
        aes_core_sbox_inst_n1623), .Y(aes_core_sbox_inst_n1407) );
  NOR4BX1 aes_core_sbox_inst_U1398 ( .AN(aes_core_sbox_inst_n1433), .B(
        aes_core_sbox_inst_n1434), .C(aes_core_sbox_inst_n277), .D(
        aes_core_sbox_inst_n1343), .Y(aes_core_sbox_inst_n1406) );
  AOI222X1 aes_core_sbox_inst_U1397 ( .A0(aes_core_sbox_inst_n184), .A1(
        aes_core_sbox_inst_n1409), .B0(aes_core_sbox_inst_n1410), .B1(
        aes_core_sbox_inst_n180), .C0(aes_core_sbox_inst_n293), .C1(
        aes_core_sbox_inst_n1411), .Y(aes_core_sbox_inst_n1408) );
  OAI222X1 aes_core_sbox_inst_U1396 ( .A0(aes_core_sbox_inst_n1406), .A1(
        aes_core_sbox_inst_n1619), .B0(aes_core_n17), .B1(
        aes_core_sbox_inst_n1407), .C0(aes_core_sbox_inst_n1408), .C1(
        aes_core_sbox_inst_n1618), .Y(aes_core_new_sboxw[13]) );
  AOI22X1 aes_core_sbox_inst_U1395 ( .A0(aes_core_sbox_inst_n56), .A1(
        aes_core_sbox_inst_n500), .B0(aes_core_sbox_inst_n501), .B1(
        aes_core_sbox_inst_n1685), .Y(aes_core_sbox_inst_n492) );
  NOR4BBX1 aes_core_sbox_inst_U1394 ( .AN(aes_core_sbox_inst_n519), .BN(
        aes_core_sbox_inst_n520), .C(aes_core_sbox_inst_n400), .D(
        aes_core_sbox_inst_n387), .Y(aes_core_sbox_inst_n491) );
  AOI222X1 aes_core_sbox_inst_U1393 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n494), .B0(aes_core_sbox_inst_n495), .B1(
        aes_core_sbox_inst_n189), .C0(aes_core_sbox_inst_n404), .C1(
        aes_core_sbox_inst_n496), .Y(aes_core_sbox_inst_n493) );
  OAI222X1 aes_core_sbox_inst_U1392 ( .A0(aes_core_sbox_inst_n491), .A1(
        aes_core_sbox_inst_n1681), .B0(aes_core_n9), .B1(
        aes_core_sbox_inst_n492), .C0(aes_core_sbox_inst_n493), .C1(
        aes_core_sbox_inst_n1680), .Y(aes_core_new_sboxw[5]) );
  INVX1 aes_core_sbox_inst_U1391 ( .A(aes_core_n6), .Y(
        aes_core_sbox_inst_n1713) );
  INVX1 aes_core_sbox_inst_U1390 ( .A(aes_core_sbox_inst_n61), .Y(
        aes_core_sbox_inst_n1595) );
  INVX1 aes_core_sbox_inst_U1389 ( .A(aes_core_n5), .Y(
        aes_core_sbox_inst_n1728) );
  BUFX3 aes_core_sbox_inst_U1388 ( .A(aes_core_sbox_inst_n1728), .Y(
        aes_core_sbox_inst_n50) );
  AOI211X1 aes_core_sbox_inst_U1387 ( .A0(aes_core_sbox_inst_n969), .A1(
        aes_core_sbox_inst_n970), .B0(aes_core_sbox_inst_n971), .C0(
        aes_core_sbox_inst_n972), .Y(aes_core_sbox_inst_n968) );
  INVX1 aes_core_sbox_inst_U1386 ( .A(aes_core_sbox_inst_n673), .Y(
        aes_core_sbox_inst_n210) );
  NOR2X1 aes_core_sbox_inst_U1385 ( .A(aes_core_sbox_inst_n209), .B(
        aes_core_sbox_inst_n206), .Y(aes_core_sbox_inst_n832) );
  INVX1 aes_core_sbox_inst_U1384 ( .A(aes_core_sbox_inst_n183), .Y(
        aes_core_sbox_inst_n182) );
  INVX1 aes_core_sbox_inst_U1383 ( .A(aes_core_sbox_inst_n440), .Y(
        aes_core_sbox_inst_n1686) );
  INVX1 aes_core_sbox_inst_U1382 ( .A(aes_core_sbox_inst_n1035), .Y(
        aes_core_sbox_inst_n1568) );
  INVX1 aes_core_sbox_inst_U1381 ( .A(aes_core_sbox_inst_n1374), .Y(
        aes_core_sbox_inst_n1624) );
  NAND3X1 aes_core_sbox_inst_U1380 ( .A(aes_core_sbox_inst_n151), .B(
        aes_core_sbox_inst_n227), .C(aes_core_sbox_inst_n637), .Y(
        aes_core_sbox_inst_n837) );
  AOI22X1 aes_core_sbox_inst_U1379 ( .A0(aes_core_sbox_inst_n81), .A1(
        aes_core_sbox_inst_n82), .B0(aes_core_sbox_inst_n85), .B1(
        aes_core_sbox_inst_n144), .Y(aes_core_sbox_inst_n1459) );
  NAND3X1 aes_core_sbox_inst_U1378 ( .A(aes_core_sbox_inst_n117), .B(
        aes_core_sbox_inst_n14), .C(aes_core_sbox_inst_n637), .Y(
        aes_core_sbox_inst_n900) );
  AOI22X1 aes_core_sbox_inst_U1377 ( .A0(aes_core_sbox_inst_n368), .A1(
        aes_core_sbox_inst_n37), .B0(aes_core_sbox_inst_n89), .B1(
        aes_core_sbox_inst_n84), .Y(aes_core_sbox_inst_n1376) );
  NOR2X1 aes_core_sbox_inst_U1376 ( .A(aes_core_sbox_inst_n1685), .B(
        aes_core_sbox_inst_n1682), .Y(aes_core_sbox_inst_n565) );
  NOR2X1 aes_core_sbox_inst_U1375 ( .A(aes_core_sbox_inst_n1567), .B(
        aes_core_sbox_inst_n450), .Y(aes_core_sbox_inst_n1190) );
  NAND2X1 aes_core_sbox_inst_U1374 ( .A(aes_core_sbox_inst_n111), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n785) );
  OAI22X1 aes_core_sbox_inst_U1373 ( .A0(aes_core_sbox_inst_n50), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n191), .B1(
        aes_core_sbox_inst_n1703), .Y(aes_core_sbox_inst_n562) );
  OAI22X1 aes_core_sbox_inst_U1372 ( .A0(aes_core_sbox_inst_n25), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n169), .B1(
        aes_core_sbox_inst_n22), .Y(aes_core_sbox_inst_n1157) );
  OAI22X1 aes_core_sbox_inst_U1371 ( .A0(aes_core_sbox_inst_n17), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n151), .B1(
        aes_core_sbox_inst_n14), .Y(aes_core_sbox_inst_n829) );
  AOI32X1 aes_core_sbox_inst_U1370 ( .A0(aes_core_sbox_inst_n33), .A1(
        aes_core_sbox_inst_n39), .A2(aes_core_sbox_inst_n79), .B0(
        aes_core_sbox_inst_n344), .B1(aes_core_sbox_inst_n80), .Y(
        aes_core_sbox_inst_n1529) );
  NOR2X1 aes_core_sbox_inst_U1369 ( .A(aes_core_sbox_inst_n18), .B(
        aes_core_sbox_inst_n17), .Y(aes_core_sbox_inst_n682) );
  NOR2X1 aes_core_sbox_inst_U1368 ( .A(aes_core_sbox_inst_n209), .B(
        aes_core_sbox_inst_n146), .Y(aes_core_sbox_inst_n859) );
  INVX1 aes_core_sbox_inst_U1367 ( .A(aes_core_sbox_inst_n155), .Y(
        aes_core_sbox_inst_n154) );
  BUFX3 aes_core_sbox_inst_U1366 ( .A(aes_core_sbox_inst_n255), .Y(
        aes_core_sbox_inst_n18) );
  INVX1 aes_core_sbox_inst_U1365 ( .A(aes_core_sbox_inst_n80), .Y(
        aes_core_sbox_inst_n1677) );
  INVX1 aes_core_sbox_inst_U1364 ( .A(aes_core_sbox_inst_n637), .Y(
        aes_core_sbox_inst_n220) );
  BUFX3 aes_core_sbox_inst_U1363 ( .A(aes_core_sbox_inst_n220), .Y(
        aes_core_sbox_inst_n13) );
  AOI2BB2X1 aes_core_sbox_inst_U1362 ( .B0(aes_core_sbox_inst_n44), .B1(
        aes_core_sbox_inst_n38), .A0N(aes_core_sbox_inst_n1645), .A1N(
        aes_core_sbox_inst_n1404), .Y(aes_core_sbox_inst_n1402) );
  AOI21X1 aes_core_sbox_inst_U1361 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n10), .B0(aes_core_sbox_inst_n358), .Y(
        aes_core_sbox_inst_n1490) );
  AOI21X1 aes_core_sbox_inst_U1360 ( .A0(aes_core_sbox_inst_n345), .A1(
        aes_core_sbox_inst_n84), .B0(aes_core_sbox_inst_n1528), .Y(
        aes_core_sbox_inst_n1526) );
  AOI222X1 aes_core_sbox_inst_U1359 ( .A0(aes_core_sbox_inst_n108), .A1(
        aes_core_sbox_inst_n119), .B0(aes_core_sbox_inst_n643), .B1(
        aes_core_sbox_inst_n159), .C0(aes_core_sbox_inst_n112), .C1(
        aes_core_sbox_inst_n136), .Y(aes_core_sbox_inst_n641) );
  NOR2BX1 aes_core_sbox_inst_U1358 ( .AN(aes_core_sbox_inst_n644), .B(
        aes_core_sbox_inst_n114), .Y(aes_core_sbox_inst_n640) );
  NAND4X1 aes_core_sbox_inst_U1357 ( .A(aes_core_sbox_inst_n639), .B(
        aes_core_sbox_inst_n224), .C(aes_core_sbox_inst_n640), .D(
        aes_core_sbox_inst_n641), .Y(aes_core_sbox_inst_n608) );
  AOI21X1 aes_core_sbox_inst_U1356 ( .A0(aes_core_sbox_inst_n36), .A1(
        aes_core_sbox_inst_n1654), .B0(aes_core_sbox_inst_n47), .Y(
        aes_core_sbox_inst_n303) );
  AOI221X1 aes_core_sbox_inst_U1355 ( .A0(aes_core_sbox_inst_n79), .A1(
        aes_core_sbox_inst_n90), .B0(aes_core_sbox_inst_n81), .B1(
        aes_core_sbox_inst_n283), .C0(aes_core_sbox_inst_n303), .Y(
        aes_core_sbox_inst_n301) );
  AOI222X1 aes_core_sbox_inst_U1354 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n82), .B0(aes_core_sbox_inst_n83), .B1(
        aes_core_sbox_inst_n47), .C0(aes_core_sbox_inst_n88), .C1(
        aes_core_sbox_inst_n45), .Y(aes_core_sbox_inst_n300) );
  AOI21X1 aes_core_sbox_inst_U1353 ( .A0(aes_core_sbox_inst_n300), .A1(
        aes_core_sbox_inst_n301), .B0(aes_core_sbox_inst_n1622), .Y(
        aes_core_sbox_inst_n299) );
  INVX1 aes_core_sbox_inst_U1352 ( .A(aes_core_sbox_inst_n1363), .Y(
        aes_core_sbox_inst_n1659) );
  AOI21X1 aes_core_sbox_inst_U1351 ( .A0(aes_core_sbox_inst_n40), .A1(
        aes_core_sbox_inst_n34), .B0(aes_core_sbox_inst_n38), .Y(
        aes_core_sbox_inst_n1405) );
  AOI22X1 aes_core_sbox_inst_U1350 ( .A0(aes_core_sbox_inst_n10), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n86), .B1(
        aes_core_sbox_inst_n40), .Y(aes_core_sbox_inst_n310) );
  NAND2BX1 aes_core_sbox_inst_U1349 ( .AN(aes_core_sbox_inst_n463), .B(
        aes_core_sbox_inst_n127), .Y(aes_core_sbox_inst_n471) );
  NAND2BX1 aes_core_sbox_inst_U1348 ( .AN(aes_core_sbox_inst_n1058), .B(
        aes_core_sbox_inst_n122), .Y(aes_core_sbox_inst_n1066) );
  NAND2BX1 aes_core_sbox_inst_U1347 ( .AN(aes_core_sbox_inst_n696), .B(
        aes_core_sbox_inst_n118), .Y(aes_core_sbox_inst_n704) );
  NAND2X1 aes_core_sbox_inst_U1346 ( .A(aes_core_sbox_inst_n410), .B(
        aes_core_sbox_inst_n5), .Y(aes_core_sbox_inst_n499) );
  NAND2X1 aes_core_sbox_inst_U1345 ( .A(aes_core_sbox_inst_n1005), .B(
        aes_core_sbox_inst_n4), .Y(aes_core_sbox_inst_n1094) );
  NAND2X1 aes_core_sbox_inst_U1344 ( .A(aes_core_sbox_inst_n643), .B(
        aes_core_sbox_inst_n9), .Y(aes_core_sbox_inst_n766) );
  OAI2BB2X1 aes_core_sbox_inst_U1343 ( .B0(aes_core_sbox_inst_n138), .B1(
        aes_core_sbox_inst_n1700), .A0N(aes_core_sbox_inst_n128), .A1N(
        aes_core_sbox_inst_n538), .Y(aes_core_sbox_inst_n543) );
  OAI2BB2X1 aes_core_sbox_inst_U1342 ( .B0(aes_core_sbox_inst_n129), .B1(
        aes_core_sbox_inst_n1582), .A0N(aes_core_sbox_inst_n123), .A1N(
        aes_core_sbox_inst_n1133), .Y(aes_core_sbox_inst_n1138) );
  OAI2BB2X1 aes_core_sbox_inst_U1341 ( .B0(aes_core_sbox_inst_n134), .B1(
        aes_core_sbox_inst_n11), .A0N(aes_core_sbox_inst_n119), .A1N(
        aes_core_sbox_inst_n805), .Y(aes_core_sbox_inst_n810) );
  AOI21X1 aes_core_sbox_inst_U1340 ( .A0(aes_core_sbox_inst_n683), .A1(
        aes_core_sbox_inst_n118), .B0(aes_core_sbox_inst_n680), .Y(
        aes_core_sbox_inst_n949) );
  AOI21X1 aes_core_sbox_inst_U1339 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n124), .B0(aes_core_sbox_inst_n1398), .Y(
        aes_core_sbox_inst_n1521) );
  AOI21X1 aes_core_sbox_inst_U1338 ( .A0(aes_core_sbox_inst_n1397), .A1(
        aes_core_sbox_inst_n80), .B0(aes_core_sbox_inst_n1368), .Y(
        aes_core_sbox_inst_n1499) );
  INVX1 aes_core_sbox_inst_U1337 ( .A(aes_core_sbox_inst_n1455), .Y(
        aes_core_sbox_inst_n1666) );
  NAND3X1 aes_core_sbox_inst_U1336 ( .A(aes_core_sbox_inst_n191), .B(
        aes_core_sbox_inst_n1704), .C(aes_core_sbox_inst_n404), .Y(
        aes_core_sbox_inst_n570) );
  NAND3X1 aes_core_sbox_inst_U1335 ( .A(aes_core_sbox_inst_n169), .B(
        aes_core_sbox_inst_n1586), .C(aes_core_sbox_inst_n999), .Y(
        aes_core_sbox_inst_n1195) );
  AOI22X1 aes_core_sbox_inst_U1334 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n199), .B0(aes_core_sbox_inst_n78), .B1(
        aes_core_sbox_inst_n138), .Y(aes_core_sbox_inst_n586) );
  AOI22X1 aes_core_sbox_inst_U1333 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n174), .B0(aes_core_sbox_inst_n104), .B1(
        aes_core_sbox_inst_n129), .Y(aes_core_sbox_inst_n1211) );
  AOI22X1 aes_core_sbox_inst_U1332 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n159), .B0(aes_core_sbox_inst_n116), .B1(
        aes_core_sbox_inst_n134), .Y(aes_core_sbox_inst_n853) );
  AOI22X1 aes_core_sbox_inst_U1331 ( .A0(aes_core_sbox_inst_n78), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n72), .B1(
        aes_core_sbox_inst_n126), .Y(aes_core_sbox_inst_n1187) );
  AOI22X1 aes_core_sbox_inst_U1330 ( .A0(aes_core_sbox_inst_n104), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n98), .B1(
        aes_core_sbox_inst_n121), .Y(aes_core_sbox_inst_n1291) );
  AOI22X1 aes_core_sbox_inst_U1329 ( .A0(aes_core_sbox_inst_n116), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n630), .B1(
        aes_core_sbox_inst_n117), .Y(aes_core_sbox_inst_n933) );
  NAND2X1 aes_core_sbox_inst_U1328 ( .A(aes_core_sbox_inst_n345), .B(
        aes_core_sbox_inst_n142), .Y(aes_core_sbox_inst_n1447) );
  AOI22X1 aes_core_sbox_inst_U1327 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n52), .B0(aes_core_sbox_inst_n71), .B1(
        aes_core_sbox_inst_n140), .Y(aes_core_sbox_inst_n549) );
  AOI22X1 aes_core_sbox_inst_U1326 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n28), .B0(aes_core_sbox_inst_n97), .B1(
        aes_core_sbox_inst_n133), .Y(aes_core_sbox_inst_n1144) );
  AOI22X1 aes_core_sbox_inst_U1325 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n19), .B0(aes_core_sbox_inst_n110), .B1(
        aes_core_sbox_inst_n136), .Y(aes_core_sbox_inst_n816) );
  AOI22X1 aes_core_sbox_inst_U1324 ( .A0(aes_core_sbox_inst_n71), .A1(
        aes_core_sbox_inst_n127), .B0(aes_core_sbox_inst_n199), .B1(
        aes_core_sbox_inst_n65), .Y(aes_core_sbox_inst_n1185) );
  AOI22X1 aes_core_sbox_inst_U1323 ( .A0(aes_core_sbox_inst_n97), .A1(
        aes_core_sbox_inst_n122), .B0(aes_core_sbox_inst_n174), .B1(
        aes_core_sbox_inst_n91), .Y(aes_core_sbox_inst_n1289) );
  AOI22X1 aes_core_sbox_inst_U1322 ( .A0(aes_core_sbox_inst_n110), .A1(
        aes_core_sbox_inst_n118), .B0(aes_core_sbox_inst_n159), .B1(
        aes_core_sbox_inst_n105), .Y(aes_core_sbox_inst_n931) );
  AOI22X1 aes_core_sbox_inst_U1321 ( .A0(aes_core_sbox_inst_n66), .A1(
        aes_core_sbox_inst_n200), .B0(aes_core_sbox_inst_n73), .B1(
        aes_core_sbox_inst_n126), .Y(aes_core_sbox_inst_n1186) );
  AOI22X1 aes_core_sbox_inst_U1320 ( .A0(aes_core_sbox_inst_n92), .A1(
        aes_core_sbox_inst_n176), .B0(aes_core_sbox_inst_n99), .B1(
        aes_core_sbox_inst_n121), .Y(aes_core_sbox_inst_n1290) );
  AOI22X1 aes_core_sbox_inst_U1319 ( .A0(aes_core_sbox_inst_n106), .A1(
        aes_core_sbox_inst_n161), .B0(aes_core_sbox_inst_n111), .B1(
        aes_core_sbox_inst_n117), .Y(aes_core_sbox_inst_n932) );
  NAND3X1 aes_core_sbox_inst_U1318 ( .A(aes_core_sbox_inst_n126), .B(
        aes_core_sbox_inst_n1703), .C(aes_core_sbox_inst_n404), .Y(
        aes_core_sbox_inst_n753) );
  NAND3X1 aes_core_sbox_inst_U1317 ( .A(aes_core_sbox_inst_n121), .B(
        aes_core_sbox_inst_n22), .C(aes_core_sbox_inst_n999), .Y(
        aes_core_sbox_inst_n1258) );
  AOI222X1 aes_core_sbox_inst_U1316 ( .A0(aes_core_sbox_inst_n1404), .A1(
        aes_core_sbox_inst_n85), .B0(aes_core_sbox_inst_n367), .B1(
        aes_core_sbox_inst_n47), .C0(aes_core_sbox_inst_n80), .C1(
        aes_core_sbox_inst_n276), .Y(aes_core_sbox_inst_n1495) );
  OAI211X1 aes_core_sbox_inst_U1315 ( .A0(aes_core_sbox_inst_n39), .A1(
        aes_core_sbox_inst_n1677), .B0(aes_core_sbox_inst_n1496), .C0(
        aes_core_sbox_inst_n1497), .Y(aes_core_sbox_inst_n1493) );
  NAND4X1 aes_core_sbox_inst_U1314 ( .A(aes_core_sbox_inst_n1447), .B(
        aes_core_sbox_inst_n1645), .C(aes_core_sbox_inst_n1391), .D(
        aes_core_sbox_inst_n1495), .Y(aes_core_sbox_inst_n1494) );
  AOI22X1 aes_core_sbox_inst_U1313 ( .A0(aes_core_sbox_inst_n263), .A1(
        aes_core_sbox_inst_n1493), .B0(aes_core_sbox_inst_n265), .B1(
        aes_core_sbox_inst_n1494), .Y(aes_core_sbox_inst_n1485) );
  NAND3X1 aes_core_sbox_inst_U1312 ( .A(aes_core_sbox_inst_n33), .B(
        aes_core_sbox_inst_n41), .C(aes_core_sbox_inst_n293), .Y(
        aes_core_sbox_inst_n1530) );
  AOI21X1 aes_core_sbox_inst_U1311 ( .A0(aes_core_sbox_inst_n463), .A1(
        aes_core_sbox_inst_n1704), .B0(aes_core_sbox_inst_n743), .Y(
        aes_core_sbox_inst_n1564) );
  AOI21X1 aes_core_sbox_inst_U1310 ( .A0(aes_core_sbox_inst_n1058), .A1(
        aes_core_sbox_inst_n1586), .B0(aes_core_sbox_inst_n1248), .Y(
        aes_core_sbox_inst_n1322) );
  AOI21X1 aes_core_sbox_inst_U1309 ( .A0(aes_core_sbox_inst_n696), .A1(
        aes_core_sbox_inst_n227), .B0(aes_core_sbox_inst_n890), .Y(
        aes_core_sbox_inst_n964) );
  AOI22X1 aes_core_sbox_inst_U1308 ( .A0(aes_core_sbox_inst_n291), .A1(
        aes_core_sbox_inst_n40), .B0(aes_core_sbox_inst_n292), .B1(
        aes_core_sbox_inst_n79), .Y(aes_core_sbox_inst_n285) );
  NAND2X1 aes_core_sbox_inst_U1307 ( .A(aes_core_sbox_inst_n67), .B(
        aes_core_sbox_inst_n66), .Y(aes_core_sbox_inst_n429) );
  NAND2X1 aes_core_sbox_inst_U1306 ( .A(aes_core_sbox_inst_n93), .B(
        aes_core_sbox_inst_n92), .Y(aes_core_sbox_inst_n1024) );
  NAND2X1 aes_core_sbox_inst_U1305 ( .A(aes_core_sbox_inst_n107), .B(
        aes_core_sbox_inst_n106), .Y(aes_core_sbox_inst_n662) );
  NAND2X1 aes_core_sbox_inst_U1304 ( .A(aes_core_sbox_inst_n79), .B(
        aes_core_sbox_inst_n321), .Y(aes_core_sbox_inst_n1362) );
  NAND2X1 aes_core_sbox_inst_U1303 ( .A(aes_core_sbox_inst_n69), .B(
        aes_core_sbox_inst_n71), .Y(aes_core_sbox_inst_n419) );
  NAND2X1 aes_core_sbox_inst_U1302 ( .A(aes_core_sbox_inst_n95), .B(
        aes_core_sbox_inst_n97), .Y(aes_core_sbox_inst_n1014) );
  NAND2X1 aes_core_sbox_inst_U1301 ( .A(aes_core_sbox_inst_n670), .B(
        aes_core_sbox_inst_n110), .Y(aes_core_sbox_inst_n652) );
  NAND3X1 aes_core_sbox_inst_U1300 ( .A(aes_core_sbox_inst_n1066), .B(
        aes_core_sbox_inst_n166), .C(aes_core_sbox_inst_n97), .Y(
        aes_core_sbox_inst_n1206) );
  NAND3X1 aes_core_sbox_inst_U1299 ( .A(aes_core_sbox_inst_n704), .B(
        aes_core_sbox_inst_n150), .C(aes_core_sbox_inst_n110), .Y(
        aes_core_sbox_inst_n848) );
  NAND3X1 aes_core_sbox_inst_U1298 ( .A(aes_core_sbox_inst_n1395), .B(
        aes_core_sbox_inst_n185), .C(aes_core_sbox_inst_n85), .Y(
        aes_core_sbox_inst_n1484) );
  AOI22X1 aes_core_sbox_inst_U1297 ( .A0(aes_core_sbox_inst_n293), .A1(
        aes_core_sbox_inst_n294), .B0(aes_core_sbox_inst_n85), .B1(
        aes_core_sbox_inst_n296), .Y(aes_core_sbox_inst_n284) );
  OAI22X1 aes_core_sbox_inst_U1296 ( .A0(aes_core_sbox_inst_n1645), .A1(
        aes_core_sbox_inst_n46), .B0(aes_core_sbox_inst_n84), .B1(
        aes_core_sbox_inst_n37), .Y(aes_core_sbox_inst_n322) );
  NAND2X1 aes_core_sbox_inst_U1295 ( .A(aes_core_sbox_inst_n73), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n518) );
  NAND2X1 aes_core_sbox_inst_U1294 ( .A(aes_core_sbox_inst_n99), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1113) );
  AOI31X1 aes_core_sbox_inst_U1293 ( .A0(aes_core_sbox_inst_n1678), .A1(
        aes_core_sbox_inst_n34), .A2(aes_core_sbox_inst_n1334), .B0(
        aes_core_sbox_inst_n1498), .Y(aes_core_sbox_inst_n1496) );
  INVX1 aes_core_sbox_inst_U1292 ( .A(aes_core_sbox_inst_n311), .Y(
        aes_core_sbox_inst_n1644) );
  AOI21X1 aes_core_sbox_inst_U1291 ( .A0(aes_core_sbox_inst_n82), .A1(
        aes_core_sbox_inst_n1673), .B0(aes_core_sbox_inst_n1644), .Y(
        aes_core_sbox_inst_n1392) );
  INVX1 aes_core_sbox_inst_U1290 ( .A(aes_core_sbox_inst_n358), .Y(
        aes_core_sbox_inst_n1667) );
  AOI31X1 aes_core_sbox_inst_U1289 ( .A0(aes_core_sbox_inst_n1391), .A1(
        aes_core_sbox_inst_n1667), .A2(aes_core_sbox_inst_n1392), .B0(
        aes_core_sbox_inst_n1622), .Y(aes_core_sbox_inst_n1390) );
  AOI22X1 aes_core_sbox_inst_U1288 ( .A0(aes_core_sbox_inst_n87), .A1(
        aes_core_sbox_inst_n79), .B0(aes_core_sbox_inst_n42), .B1(
        aes_core_sbox_inst_n86), .Y(aes_core_sbox_inst_n342) );
  AOI21X1 aes_core_sbox_inst_U1287 ( .A0(aes_core_sbox_inst_n142), .A1(
        aes_core_sbox_inst_n86), .B0(aes_core_sbox_inst_n1387), .Y(
        aes_core_sbox_inst_n1445) );
  AOI32X1 aes_core_sbox_inst_U1286 ( .A0(aes_core_sbox_inst_n125), .A1(
        aes_core_sbox_inst_n39), .A2(aes_core_sbox_inst_n1446), .B0(
        aes_core_sbox_inst_n79), .B1(aes_core_sbox_inst_n272), .Y(
        aes_core_sbox_inst_n1444) );
  OAI211X1 aes_core_sbox_inst_U1285 ( .A0(aes_core_sbox_inst_n1660), .A1(
        aes_core_sbox_inst_n1677), .B0(aes_core_sbox_inst_n1444), .C0(
        aes_core_sbox_inst_n1445), .Y(aes_core_sbox_inst_n1443) );
  AOI222X1 aes_core_sbox_inst_U1284 ( .A0(aes_core_sbox_inst_n116), .A1(
        aes_core_sbox_inst_n20), .B0(aes_core_sbox_inst_n643), .B1(
        aes_core_sbox_inst_n136), .C0(aes_core_sbox_inst_n112), .C1(
        aes_core_sbox_inst_n9), .Y(aes_core_sbox_inst_n666) );
  AOI31X1 aes_core_sbox_inst_U1283 ( .A0(aes_core_sbox_inst_n664), .A1(
        aes_core_sbox_inst_n665), .A2(aes_core_sbox_inst_n666), .B0(
        aes_core_sbox_inst_n149), .Y(aes_core_sbox_inst_n660) );
  NOR2X1 aes_core_sbox_inst_U1282 ( .A(aes_core_sbox_inst_n82), .B(
        aes_core_sbox_inst_n321), .Y(aes_core_sbox_inst_n1446) );
  NOR2X1 aes_core_sbox_inst_U1281 ( .A(aes_core_sbox_inst_n79), .B(
        aes_core_sbox_inst_n179), .Y(aes_core_sbox_inst_n1344) );
  AOI31X1 aes_core_sbox_inst_U1280 ( .A0(aes_core_sbox_inst_n769), .A1(
        aes_core_sbox_inst_n802), .A2(aes_core_sbox_inst_n650), .B0(
        aes_core_sbox_inst_n148), .Y(aes_core_sbox_inst_n929) );
  AOI31X1 aes_core_sbox_inst_U1279 ( .A0(aes_core_sbox_inst_n933), .A1(
        aes_core_sbox_inst_n709), .A2(aes_core_sbox_inst_n934), .B0(
        aes_core_sbox_inst_n147), .Y(aes_core_sbox_inst_n928) );
  AOI21X1 aes_core_sbox_inst_U1278 ( .A0(aes_core_sbox_inst_n931), .A1(
        aes_core_sbox_inst_n932), .B0(aes_core_sbox_inst_n215), .Y(
        aes_core_sbox_inst_n930) );
  OAI31X1 aes_core_sbox_inst_U1277 ( .A0(aes_core_sbox_inst_n928), .A1(
        aes_core_sbox_inst_n929), .A2(aes_core_sbox_inst_n930), .B0(
        aes_core_sbox_inst_n209), .Y(aes_core_sbox_inst_n919) );
  NOR2X1 aes_core_sbox_inst_U1276 ( .A(aes_core_sbox_inst_n73), .B(
        aes_core_sbox_inst_n66), .Y(aes_core_sbox_inst_n385) );
  NOR2X1 aes_core_sbox_inst_U1275 ( .A(aes_core_sbox_inst_n99), .B(
        aes_core_sbox_inst_n92), .Y(aes_core_sbox_inst_n980) );
  NOR2X1 aes_core_sbox_inst_U1274 ( .A(aes_core_sbox_inst_n111), .B(
        aes_core_sbox_inst_n106), .Y(aes_core_sbox_inst_n618) );
  NAND2X1 aes_core_sbox_inst_U1273 ( .A(aes_core_sbox_inst_n3), .B(
        aes_core_sbox_inst_n138), .Y(aes_core_sbox_inst_n553) );
  NAND2X1 aes_core_sbox_inst_U1272 ( .A(aes_core_sbox_inst_n1045), .B(
        aes_core_sbox_inst_n129), .Y(aes_core_sbox_inst_n1148) );
  NAND2X1 aes_core_sbox_inst_U1271 ( .A(aes_core_sbox_inst_n683), .B(
        aes_core_sbox_inst_n134), .Y(aes_core_sbox_inst_n820) );
  AOI221X1 aes_core_sbox_inst_U1270 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n1545), .B0(aes_core_sbox_inst_n6), .B1(
        aes_core_sbox_inst_n75), .C0(aes_core_sbox_inst_n576), .Y(
        aes_core_sbox_inst_n1538) );
  AOI221X1 aes_core_sbox_inst_U1269 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n1303), .B0(aes_core_sbox_inst_n7), .B1(
        aes_core_sbox_inst_n101), .C0(aes_core_sbox_inst_n1201), .Y(
        aes_core_sbox_inst_n1296) );
  AOI221X1 aes_core_sbox_inst_U1268 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n945), .B0(aes_core_sbox_inst_n8), .B1(
        aes_core_sbox_inst_n113), .C0(aes_core_sbox_inst_n843), .Y(
        aes_core_sbox_inst_n938) );
  AOI32X1 aes_core_sbox_inst_U1267 ( .A0(aes_core_sbox_inst_n1703), .A1(
        aes_core_sbox_inst_n1732), .A2(aes_core_sbox_inst_n67), .B0(
        aes_core_sbox_inst_n561), .B1(aes_core_sbox_inst_n5), .Y(
        aes_core_sbox_inst_n748) );
  AOI32X1 aes_core_sbox_inst_U1266 ( .A0(aes_core_sbox_inst_n22), .A1(
        aes_core_sbox_inst_n27), .A2(aes_core_sbox_inst_n93), .B0(
        aes_core_sbox_inst_n1156), .B1(aes_core_sbox_inst_n4), .Y(
        aes_core_sbox_inst_n1253) );
  AOI32X1 aes_core_sbox_inst_U1265 ( .A0(aes_core_sbox_inst_n14), .A1(
        aes_core_sbox_inst_n18), .A2(aes_core_sbox_inst_n107), .B0(
        aes_core_sbox_inst_n828), .B1(aes_core_sbox_inst_n9), .Y(
        aes_core_sbox_inst_n895) );
  NAND2X1 aes_core_sbox_inst_U1264 ( .A(aes_core_sbox_inst_n1651), .B(
        aes_core_sbox_inst_n1660), .Y(aes_core_sbox_inst_n1386) );
  AOI222X1 aes_core_sbox_inst_U1263 ( .A0(aes_core_sbox_inst_n81), .A1(
        aes_core_sbox_inst_n272), .B0(aes_core_sbox_inst_n1386), .B1(
        aes_core_sbox_inst_n47), .C0(aes_core_sbox_inst_n80), .C1(
        aes_core_sbox_inst_n275), .Y(aes_core_sbox_inst_n1385) );
  AOI222X1 aes_core_sbox_inst_U1262 ( .A0(aes_core_sbox_inst_n87), .A1(
        aes_core_sbox_inst_n1673), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n86), .C0(aes_core_sbox_inst_n84), .C1(
        aes_core_sbox_inst_n82), .Y(aes_core_sbox_inst_n1384) );
  OAI221X1 aes_core_sbox_inst_U1261 ( .A0(aes_core_sbox_inst_n35), .A1(
        aes_core_sbox_inst_n336), .B0(aes_core_sbox_inst_n1677), .B1(
        aes_core_sbox_inst_n1651), .C0(aes_core_sbox_inst_n337), .Y(
        aes_core_sbox_inst_n335) );
  AOI222X1 aes_core_sbox_inst_U1260 ( .A0(aes_core_sbox_inst_n69), .A1(
        aes_core_sbox_inst_n66), .B0(aes_core_sbox_inst_n561), .B1(
        aes_core_sbox_inst_n67), .C0(aes_core_sbox_inst_n78), .C1(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n559) );
  AOI222X1 aes_core_sbox_inst_U1259 ( .A0(aes_core_sbox_inst_n95), .A1(
        aes_core_sbox_inst_n92), .B0(aes_core_sbox_inst_n1156), .B1(
        aes_core_sbox_inst_n93), .C0(aes_core_sbox_inst_n104), .C1(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1154) );
  AOI222X1 aes_core_sbox_inst_U1258 ( .A0(aes_core_sbox_inst_n670), .A1(
        aes_core_sbox_inst_n106), .B0(aes_core_sbox_inst_n828), .B1(
        aes_core_sbox_inst_n107), .C0(aes_core_sbox_inst_n116), .C1(
        aes_core_sbox_inst_n160), .Y(aes_core_sbox_inst_n826) );
  AOI211X1 aes_core_sbox_inst_U1257 ( .A0(aes_core_sbox_inst_n446), .A1(
        aes_core_sbox_inst_n200), .B0(aes_core_sbox_inst_n447), .C0(
        aes_core_sbox_inst_n448), .Y(aes_core_sbox_inst_n445) );
  AOI211X1 aes_core_sbox_inst_U1256 ( .A0(aes_core_sbox_inst_n1041), .A1(
        aes_core_sbox_inst_n177), .B0(aes_core_sbox_inst_n1042), .C0(
        aes_core_sbox_inst_n1043), .Y(aes_core_sbox_inst_n1040) );
  AOI211X1 aes_core_sbox_inst_U1255 ( .A0(aes_core_sbox_inst_n679), .A1(
        aes_core_sbox_inst_n161), .B0(aes_core_sbox_inst_n680), .C0(
        aes_core_sbox_inst_n681), .Y(aes_core_sbox_inst_n678) );
  NOR2X1 aes_core_sbox_inst_U1254 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n50), .Y(aes_core_sbox_inst_n449) );
  NOR2X1 aes_core_sbox_inst_U1253 ( .A(aes_core_sbox_inst_n27), .B(
        aes_core_sbox_inst_n25), .Y(aes_core_sbox_inst_n1044) );
  NOR2X1 aes_core_sbox_inst_U1252 ( .A(aes_core_sbox_inst_n38), .B(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n1379) );
  NAND2X1 aes_core_sbox_inst_U1251 ( .A(aes_core_sbox_inst_n88), .B(
        aes_core_sbox_inst_n79), .Y(aes_core_sbox_inst_n319) );
  AOI222X1 aes_core_sbox_inst_U1250 ( .A0(aes_core_sbox_inst_n490), .A1(
        aes_core_sbox_inst_n66), .B0(aes_core_sbox_inst_n77), .B1(
        aes_core_sbox_inst_n200), .C0(aes_core_sbox_inst_n69), .C1(
        aes_core_sbox_inst_n68), .Y(aes_core_sbox_inst_n588) );
  AOI222X1 aes_core_sbox_inst_U1249 ( .A0(aes_core_sbox_inst_n1085), .A1(
        aes_core_sbox_inst_n92), .B0(aes_core_sbox_inst_n103), .B1(
        aes_core_sbox_inst_n175), .C0(aes_core_sbox_inst_n95), .C1(
        aes_core_sbox_inst_n94), .Y(aes_core_sbox_inst_n1213) );
  AOI222X1 aes_core_sbox_inst_U1248 ( .A0(aes_core_sbox_inst_n723), .A1(
        aes_core_sbox_inst_n106), .B0(aes_core_sbox_inst_n115), .B1(
        aes_core_sbox_inst_n161), .C0(aes_core_sbox_inst_n670), .C1(
        aes_core_sbox_inst_n108), .Y(aes_core_sbox_inst_n855) );
  AOI222X1 aes_core_sbox_inst_U1247 ( .A0(aes_core_sbox_inst_n1404), .A1(
        aes_core_sbox_inst_n321), .B0(aes_core_sbox_inst_n83), .B1(
        aes_core_sbox_inst_n47), .C0(aes_core_sbox_inst_n356), .C1(
        aes_core_sbox_inst_n84), .Y(aes_core_sbox_inst_n1491) );
  NOR4BX1 aes_core_sbox_inst_U1246 ( .AN(aes_core_sbox_inst_n1468), .B(
        aes_core_sbox_inst_n315), .C(aes_core_sbox_inst_n1469), .D(
        aes_core_sbox_inst_n346), .Y(aes_core_sbox_inst_n1467) );
  AOI221X1 aes_core_sbox_inst_U1245 ( .A0(aes_core_sbox_inst_n356), .A1(
        aes_core_sbox_inst_n79), .B0(aes_core_sbox_inst_n88), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n1455), .Y(
        aes_core_sbox_inst_n1465) );
  AOI211X1 aes_core_sbox_inst_U1244 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n34), .B0(aes_core_sbox_inst_n294), .C0(
        aes_core_sbox_inst_n82), .Y(aes_core_sbox_inst_n1466) );
  OAI222X1 aes_core_sbox_inst_U1243 ( .A0(aes_core_sbox_inst_n179), .A1(
        aes_core_sbox_inst_n1465), .B0(aes_core_sbox_inst_n1466), .B1(
        aes_core_sbox_inst_n31), .C0(aes_core_sbox_inst_n1467), .C1(
        aes_core_sbox_inst_n181), .Y(aes_core_sbox_inst_n1457) );
  AOI221X1 aes_core_sbox_inst_U1242 ( .A0(aes_core_sbox_inst_n85), .A1(
        aes_core_sbox_inst_n47), .B0(aes_core_sbox_inst_n321), .B1(
        aes_core_sbox_inst_n125), .C0(aes_core_sbox_inst_n333), .Y(
        aes_core_sbox_inst_n332) );
  NOR2X1 aes_core_sbox_inst_U1241 ( .A(aes_core_sbox_inst_n1697), .B(
        aes_core_sbox_inst_n50), .Y(aes_core_sbox_inst_n573) );
  NOR2X1 aes_core_sbox_inst_U1240 ( .A(aes_core_sbox_inst_n34), .B(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n315) );
  INVX1 aes_core_sbox_inst_U1239 ( .A(aes_core_sbox_inst_n1514), .Y(
        aes_core_sbox_inst_n1662) );
  AOI221X1 aes_core_sbox_inst_U1238 ( .A0(aes_core_sbox_inst_n90), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n356), .B1(
        aes_core_sbox_inst_n43), .C0(aes_core_sbox_inst_n1662), .Y(
        aes_core_sbox_inst_n1522) );
  AOI222X1 aes_core_sbox_inst_U1237 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n449), .B1(
        aes_core_sbox_inst_n126), .C0(aes_core_sbox_inst_n3), .C1(
        aes_core_sbox_inst_n192), .Y(aes_core_sbox_inst_n444) );
  AOI222X1 aes_core_sbox_inst_U1236 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n1044), .B1(
        aes_core_sbox_inst_n121), .C0(aes_core_sbox_inst_n1045), .C1(
        aes_core_sbox_inst_n170), .Y(aes_core_sbox_inst_n1039) );
  AOI222X1 aes_core_sbox_inst_U1235 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n155), .B0(aes_core_sbox_inst_n682), .B1(
        aes_core_sbox_inst_n117), .C0(aes_core_sbox_inst_n683), .C1(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n677) );
  AOI222X1 aes_core_sbox_inst_U1234 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n128), .B0(aes_core_sbox_inst_n446), .B1(
        aes_core_sbox_inst_n69), .C0(aes_core_sbox_inst_n74), .C1(
        aes_core_sbox_inst_n6), .Y(aes_core_sbox_inst_n555) );
  AOI222X1 aes_core_sbox_inst_U1233 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n123), .B0(aes_core_sbox_inst_n1041), .B1(
        aes_core_sbox_inst_n95), .C0(aes_core_sbox_inst_n100), .C1(
        aes_core_sbox_inst_n7), .Y(aes_core_sbox_inst_n1150) );
  AOI222X1 aes_core_sbox_inst_U1232 ( .A0(aes_core_sbox_inst_n356), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n84), .B1(
        aes_core_sbox_inst_n90), .C0(aes_core_sbox_inst_n83), .C1(
        aes_core_sbox_inst_n44), .Y(aes_core_sbox_inst_n355) );
  AOI222X1 aes_core_sbox_inst_U1231 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n119), .B0(aes_core_sbox_inst_n679), .B1(
        aes_core_sbox_inst_n670), .C0(aes_core_sbox_inst_n112), .C1(
        aes_core_sbox_inst_n8), .Y(aes_core_sbox_inst_n822) );
  AOI222X1 aes_core_sbox_inst_U1230 ( .A0(aes_core_sbox_inst_n71), .A1(
        aes_core_sbox_inst_n199), .B0(aes_core_sbox_inst_n545), .B1(
        aes_core_sbox_inst_n67), .C0(aes_core_sbox_inst_n74), .C1(
        aes_core_sbox_inst_n139), .Y(aes_core_sbox_inst_n1565) );
  AOI222X1 aes_core_sbox_inst_U1229 ( .A0(aes_core_sbox_inst_n97), .A1(
        aes_core_sbox_inst_n174), .B0(aes_core_sbox_inst_n1140), .B1(
        aes_core_sbox_inst_n93), .C0(aes_core_sbox_inst_n100), .C1(
        aes_core_sbox_inst_n130), .Y(aes_core_sbox_inst_n1323) );
  AOI222X1 aes_core_sbox_inst_U1228 ( .A0(aes_core_sbox_inst_n110), .A1(
        aes_core_sbox_inst_n159), .B0(aes_core_sbox_inst_n812), .B1(
        aes_core_sbox_inst_n107), .C0(aes_core_sbox_inst_n112), .C1(
        aes_core_sbox_inst_n135), .Y(aes_core_sbox_inst_n965) );
  AOI222X1 aes_core_sbox_inst_U1227 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n90), .B0(aes_core_sbox_inst_n1380), .B1(
        aes_core_sbox_inst_n84), .C0(aes_core_sbox_inst_n89), .C1(
        aes_core_sbox_inst_n45), .Y(aes_core_sbox_inst_n1464) );
  INVX1 aes_core_sbox_inst_U1226 ( .A(aes_core_sbox_inst_n488), .Y(
        aes_core_sbox_inst_n1691) );
  INVX1 aes_core_sbox_inst_U1225 ( .A(aes_core_sbox_inst_n1083), .Y(
        aes_core_sbox_inst_n1573) );
  INVX1 aes_core_sbox_inst_U1224 ( .A(aes_core_sbox_inst_n198), .Y(
        aes_core_sbox_inst_n197) );
  INVX1 aes_core_sbox_inst_U1223 ( .A(aes_core_sbox_inst_n197), .Y(
        aes_core_sbox_inst_n203) );
  INVX1 aes_core_sbox_inst_U1222 ( .A(aes_core_n18), .Y(
        aes_core_sbox_inst_n178) );
  INVX1 aes_core_sbox_inst_U1221 ( .A(aes_core_sbox_inst_n158), .Y(
        aes_core_sbox_inst_n157) );
  INVX1 aes_core_sbox_inst_U1220 ( .A(aes_core_sbox_inst_n198), .Y(
        aes_core_sbox_inst_n196) );
  INVX1 aes_core_sbox_inst_U1219 ( .A(aes_core_sbox_inst_n158), .Y(
        aes_core_sbox_inst_n156) );
  INVX1 aes_core_sbox_inst_U1218 ( .A(aes_core_sbox_inst_n321), .Y(
        aes_core_sbox_inst_n1655) );
  BUFX3 aes_core_sbox_inst_U1217 ( .A(aes_core_sbox_inst_n1655), .Y(
        aes_core_sbox_inst_n33) );
  OAI222X1 aes_core_sbox_inst_U1216 ( .A0(aes_core_sbox_inst_n184), .A1(
        aes_core_sbox_inst_n1402), .B0(aes_core_sbox_inst_n1403), .B1(
        aes_core_sbox_inst_n181), .C0(aes_core_sbox_inst_n1404), .C1(
        aes_core_sbox_inst_n37), .Y(aes_core_sbox_inst_n1401) );
  AOI21X1 aes_core_sbox_inst_U1215 ( .A0(aes_core_sbox_inst_n1671), .A1(
        aes_core_sbox_inst_n1648), .B0(aes_core_sbox_inst_n1630), .Y(
        aes_core_sbox_inst_n1400) );
  NOR2X1 aes_core_sbox_inst_U1214 ( .A(aes_core_sbox_inst_n1405), .B(
        aes_core_sbox_inst_n1636), .Y(aes_core_sbox_inst_n1399) );
  OR4X2 aes_core_sbox_inst_U1213 ( .A(aes_core_sbox_inst_n1398), .B(
        aes_core_sbox_inst_n1399), .C(aes_core_sbox_inst_n1400), .D(
        aes_core_sbox_inst_n1401), .Y(aes_core_sbox_inst_n1388) );
  OAI2BB1X1 aes_core_sbox_inst_U1212 ( .A0N(aes_core_sbox_inst_n126), .A1N(
        aes_core_sbox_inst_n74), .B0(aes_core_sbox_inst_n1717), .Y(
        aes_core_sbox_inst_n517) );
  OAI2BB1X1 aes_core_sbox_inst_U1211 ( .A0N(aes_core_sbox_inst_n121), .A1N(
        aes_core_sbox_inst_n100), .B0(aes_core_sbox_inst_n1599), .Y(
        aes_core_sbox_inst_n1112) );
  OAI2BB1X1 aes_core_sbox_inst_U1210 ( .A0N(aes_core_sbox_inst_n117), .A1N(
        aes_core_sbox_inst_n112), .B0(aes_core_sbox_inst_n240), .Y(
        aes_core_sbox_inst_n784) );
  INVX1 aes_core_sbox_inst_U1209 ( .A(aes_core_sbox_inst_n79), .Y(
        aes_core_sbox_inst_n1675) );
  INVX1 aes_core_sbox_inst_U1208 ( .A(aes_core_sbox_inst_n404), .Y(
        aes_core_sbox_inst_n1696) );
  BUFX3 aes_core_sbox_inst_U1207 ( .A(aes_core_sbox_inst_n1696), .Y(
        aes_core_sbox_inst_n48) );
  INVX1 aes_core_sbox_inst_U1206 ( .A(aes_core_sbox_inst_n999), .Y(
        aes_core_sbox_inst_n1578) );
  BUFX3 aes_core_sbox_inst_U1205 ( .A(aes_core_sbox_inst_n1578), .Y(
        aes_core_sbox_inst_n21) );
  INVX1 aes_core_sbox_inst_U1204 ( .A(aes_core_sbox_inst_n293), .Y(
        aes_core_sbox_inst_n1635) );
  BUFX3 aes_core_sbox_inst_U1203 ( .A(aes_core_sbox_inst_n1635), .Y(
        aes_core_sbox_inst_n31) );
  NOR2X1 aes_core_sbox_inst_U1202 ( .A(aes_core_sbox_inst_n80), .B(
        aes_core_sbox_inst_n79), .Y(aes_core_sbox_inst_n302) );
  BUFX3 aes_core_sbox_inst_U1201 ( .A(aes_core_sbox_inst_n302), .Y(
        aes_core_sbox_inst_n81) );
  AOI21X1 aes_core_sbox_inst_U1200 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n283), .B0(aes_core_sbox_inst_n369), .Y(
        aes_core_sbox_inst_n1519) );
  OAI211X1 aes_core_sbox_inst_U1199 ( .A0(aes_core_sbox_inst_n192), .A1(
        aes_core_sbox_inst_n1720), .B0(aes_core_sbox_inst_n416), .C0(
        aes_core_sbox_inst_n459), .Y(aes_core_sbox_inst_n454) );
  AOI22X1 aes_core_sbox_inst_U1198 ( .A0(aes_core_sbox_inst_n186), .A1(
        aes_core_sbox_inst_n454), .B0(aes_core_sbox_inst_n455), .B1(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n451) );
  AOI22X1 aes_core_sbox_inst_U1197 ( .A0(aes_core_sbox_inst_n392), .A1(
        aes_core_sbox_inst_n138), .B0(aes_core_sbox_inst_n69), .B1(
        aes_core_sbox_inst_n453), .Y(aes_core_sbox_inst_n452) );
  AOI21X1 aes_core_sbox_inst_U1196 ( .A0(aes_core_sbox_inst_n451), .A1(
        aes_core_sbox_inst_n452), .B0(aes_core_sbox_inst_n1685), .Y(
        aes_core_sbox_inst_n442) );
  OAI211X1 aes_core_sbox_inst_U1195 ( .A0(aes_core_sbox_inst_n170), .A1(
        aes_core_sbox_inst_n24), .B0(aes_core_sbox_inst_n1011), .C0(
        aes_core_sbox_inst_n1054), .Y(aes_core_sbox_inst_n1049) );
  AOI22X1 aes_core_sbox_inst_U1194 ( .A0(aes_core_sbox_inst_n164), .A1(
        aes_core_sbox_inst_n1049), .B0(aes_core_sbox_inst_n1050), .B1(
        aes_core_sbox_inst_n167), .Y(aes_core_sbox_inst_n1046) );
  AOI22X1 aes_core_sbox_inst_U1193 ( .A0(aes_core_sbox_inst_n987), .A1(
        aes_core_sbox_inst_n129), .B0(aes_core_sbox_inst_n95), .B1(
        aes_core_sbox_inst_n1048), .Y(aes_core_sbox_inst_n1047) );
  AOI21X1 aes_core_sbox_inst_U1192 ( .A0(aes_core_sbox_inst_n1046), .A1(
        aes_core_sbox_inst_n1047), .B0(aes_core_sbox_inst_n1567), .Y(
        aes_core_sbox_inst_n1037) );
  OAI211X1 aes_core_sbox_inst_U1191 ( .A0(aes_core_sbox_inst_n154), .A1(
        aes_core_sbox_inst_n243), .B0(aes_core_sbox_inst_n649), .C0(
        aes_core_sbox_inst_n692), .Y(aes_core_sbox_inst_n687) );
  AOI22X1 aes_core_sbox_inst_U1190 ( .A0(aes_core_sbox_inst_n146), .A1(
        aes_core_sbox_inst_n687), .B0(aes_core_sbox_inst_n688), .B1(
        aes_core_sbox_inst_n149), .Y(aes_core_sbox_inst_n684) );
  AOI22X1 aes_core_sbox_inst_U1189 ( .A0(aes_core_sbox_inst_n625), .A1(
        aes_core_sbox_inst_n134), .B0(aes_core_sbox_inst_n670), .B1(
        aes_core_sbox_inst_n686), .Y(aes_core_sbox_inst_n685) );
  AOI21X1 aes_core_sbox_inst_U1188 ( .A0(aes_core_sbox_inst_n684), .A1(
        aes_core_sbox_inst_n685), .B0(aes_core_sbox_inst_n209), .Y(
        aes_core_sbox_inst_n675) );
  AOI21X1 aes_core_sbox_inst_U1187 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n52), .B0(aes_core_sbox_inst_n477), .Y(
        aes_core_sbox_inst_n587) );
  AOI21X1 aes_core_sbox_inst_U1186 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n28), .B0(aes_core_sbox_inst_n1072), .Y(
        aes_core_sbox_inst_n1212) );
  AOI21X1 aes_core_sbox_inst_U1185 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n19), .B0(aes_core_sbox_inst_n710), .Y(
        aes_core_sbox_inst_n854) );
  AOI31X1 aes_core_sbox_inst_U1184 ( .A0(aes_core_sbox_inst_n200), .A1(
        aes_core_sbox_inst_n189), .A2(aes_core_sbox_inst_n75), .B0(
        aes_core_sbox_inst_n405), .Y(aes_core_sbox_inst_n1171) );
  AOI22X1 aes_core_sbox_inst_U1183 ( .A0(aes_core_sbox_inst_n453), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n573), .B1(
        aes_core_sbox_inst_n67), .Y(aes_core_sbox_inst_n1169) );
  AOI22X1 aes_core_sbox_inst_U1182 ( .A0(aes_core_sbox_inst_n404), .A1(
        aes_core_sbox_inst_n562), .B0(aes_core_sbox_inst_n71), .B1(
        aes_core_sbox_inst_n406), .Y(aes_core_sbox_inst_n1168) );
  NAND4X1 aes_core_sbox_inst_U1181 ( .A(aes_core_sbox_inst_n1168), .B(
        aes_core_sbox_inst_n1169), .C(aes_core_sbox_inst_n1170), .D(
        aes_core_sbox_inst_n1171), .Y(aes_core_sbox_inst_n1161) );
  AOI31X1 aes_core_sbox_inst_U1180 ( .A0(aes_core_sbox_inst_n175), .A1(
        aes_core_sbox_inst_n167), .A2(aes_core_sbox_inst_n101), .B0(
        aes_core_sbox_inst_n1000), .Y(aes_core_sbox_inst_n1275) );
  AOI22X1 aes_core_sbox_inst_U1179 ( .A0(aes_core_sbox_inst_n1048), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n1198), .B1(
        aes_core_sbox_inst_n93), .Y(aes_core_sbox_inst_n1273) );
  AOI22X1 aes_core_sbox_inst_U1178 ( .A0(aes_core_sbox_inst_n999), .A1(
        aes_core_sbox_inst_n1157), .B0(aes_core_sbox_inst_n97), .B1(
        aes_core_sbox_inst_n1001), .Y(aes_core_sbox_inst_n1272) );
  NAND4X1 aes_core_sbox_inst_U1177 ( .A(aes_core_sbox_inst_n1272), .B(
        aes_core_sbox_inst_n1273), .C(aes_core_sbox_inst_n1274), .D(
        aes_core_sbox_inst_n1275), .Y(aes_core_sbox_inst_n1265) );
  AOI31X1 aes_core_sbox_inst_U1176 ( .A0(aes_core_sbox_inst_n161), .A1(
        aes_core_sbox_inst_n148), .A2(aes_core_sbox_inst_n113), .B0(
        aes_core_sbox_inst_n638), .Y(aes_core_sbox_inst_n917) );
  AOI22X1 aes_core_sbox_inst_U1175 ( .A0(aes_core_sbox_inst_n637), .A1(
        aes_core_sbox_inst_n829), .B0(aes_core_sbox_inst_n110), .B1(
        aes_core_sbox_inst_n639), .Y(aes_core_sbox_inst_n914) );
  AOI22X1 aes_core_sbox_inst_U1174 ( .A0(aes_core_sbox_inst_n686), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n840), .B1(
        aes_core_sbox_inst_n107), .Y(aes_core_sbox_inst_n915) );
  NAND4X1 aes_core_sbox_inst_U1173 ( .A(aes_core_sbox_inst_n914), .B(
        aes_core_sbox_inst_n915), .C(aes_core_sbox_inst_n916), .D(
        aes_core_sbox_inst_n917), .Y(aes_core_sbox_inst_n907) );
  AOI21X1 aes_core_sbox_inst_U1172 ( .A0(aes_core_sbox_inst_n1724), .A1(
        aes_core_sbox_inst_n1706), .B0(aes_core_sbox_inst_n126), .Y(
        aes_core_sbox_inst_n498) );
  INVX1 aes_core_sbox_inst_U1171 ( .A(aes_core_sbox_inst_n499), .Y(
        aes_core_sbox_inst_n1729) );
  AOI211X1 aes_core_sbox_inst_U1170 ( .A0(aes_core_sbox_inst_n78), .A1(
        aes_core_sbox_inst_n139), .B0(aes_core_sbox_inst_n1729), .C0(
        aes_core_sbox_inst_n498), .Y(aes_core_sbox_inst_n497) );
  NAND4X1 aes_core_sbox_inst_U1169 ( .A(aes_core_sbox_inst_n419), .B(
        aes_core_sbox_inst_n395), .C(aes_core_sbox_inst_n1701), .D(
        aes_core_sbox_inst_n497), .Y(aes_core_sbox_inst_n494) );
  AOI21X1 aes_core_sbox_inst_U1168 ( .A0(aes_core_sbox_inst_n1606), .A1(
        aes_core_sbox_inst_n1588), .B0(aes_core_sbox_inst_n121), .Y(
        aes_core_sbox_inst_n1093) );
  INVX1 aes_core_sbox_inst_U1167 ( .A(aes_core_sbox_inst_n1094), .Y(
        aes_core_sbox_inst_n1611) );
  AOI211X1 aes_core_sbox_inst_U1166 ( .A0(aes_core_sbox_inst_n104), .A1(
        aes_core_sbox_inst_n130), .B0(aes_core_sbox_inst_n1611), .C0(
        aes_core_sbox_inst_n1093), .Y(aes_core_sbox_inst_n1092) );
  NAND4X1 aes_core_sbox_inst_U1165 ( .A(aes_core_sbox_inst_n1014), .B(
        aes_core_sbox_inst_n990), .C(aes_core_sbox_inst_n1583), .D(
        aes_core_sbox_inst_n1092), .Y(aes_core_sbox_inst_n1089) );
  AOI21X1 aes_core_sbox_inst_U1164 ( .A0(aes_core_sbox_inst_n247), .A1(
        aes_core_sbox_inst_n229), .B0(aes_core_sbox_inst_n117), .Y(
        aes_core_sbox_inst_n765) );
  INVX1 aes_core_sbox_inst_U1163 ( .A(aes_core_sbox_inst_n766), .Y(
        aes_core_sbox_inst_n252) );
  AOI211X1 aes_core_sbox_inst_U1162 ( .A0(aes_core_sbox_inst_n116), .A1(
        aes_core_sbox_inst_n135), .B0(aes_core_sbox_inst_n252), .C0(
        aes_core_sbox_inst_n765), .Y(aes_core_sbox_inst_n764) );
  NAND4X1 aes_core_sbox_inst_U1161 ( .A(aes_core_sbox_inst_n652), .B(
        aes_core_sbox_inst_n628), .C(aes_core_sbox_inst_n224), .D(
        aes_core_sbox_inst_n764), .Y(aes_core_sbox_inst_n761) );
  AOI21X1 aes_core_sbox_inst_U1160 ( .A0(aes_core_sbox_inst_n1661), .A1(
        aes_core_sbox_inst_n1638), .B0(aes_core_sbox_inst_n40), .Y(
        aes_core_sbox_inst_n1414) );
  AOI221X1 aes_core_sbox_inst_U1159 ( .A0(aes_core_sbox_inst_n84), .A1(
        aes_core_sbox_inst_n85), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n10), .C0(aes_core_sbox_inst_n1414), .Y(
        aes_core_sbox_inst_n1413) );
  NAND4X1 aes_core_sbox_inst_U1158 ( .A(aes_core_sbox_inst_n1650), .B(
        aes_core_sbox_inst_n1340), .C(aes_core_sbox_inst_n1412), .D(
        aes_core_sbox_inst_n1413), .Y(aes_core_sbox_inst_n1409) );
  NAND4X1 aes_core_sbox_inst_U1157 ( .A(aes_core_sbox_inst_n1340), .B(
        aes_core_sbox_inst_n36), .C(aes_core_sbox_inst_n353), .D(
        aes_core_sbox_inst_n1512), .Y(aes_core_sbox_inst_n1511) );
  AOI22X1 aes_core_sbox_inst_U1156 ( .A0(aes_core_sbox_inst_n179), .A1(
        aes_core_sbox_inst_n1510), .B0(aes_core_sbox_inst_n1511), .B1(
        aes_core_sbox_inst_n182), .Y(aes_core_sbox_inst_n1508) );
  AOI221X1 aes_core_sbox_inst_U1155 ( .A0(aes_core_sbox_inst_n307), .A1(
        aes_core_sbox_inst_n125), .B0(aes_core_sbox_inst_n290), .B1(
        aes_core_sbox_inst_n81), .C0(aes_core_sbox_inst_n1358), .Y(
        aes_core_sbox_inst_n1509) );
  AOI21X1 aes_core_sbox_inst_U1154 ( .A0(aes_core_sbox_inst_n1508), .A1(
        aes_core_sbox_inst_n1509), .B0(aes_core_sbox_inst_n1618), .Y(
        aes_core_sbox_inst_n1507) );
  AOI222X1 aes_core_sbox_inst_U1153 ( .A0(aes_core_sbox_inst_n65), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n75), .B1(
        aes_core_sbox_inst_n70), .C0(aes_core_sbox_inst_n72), .C1(
        aes_core_sbox_inst_n53), .Y(aes_core_sbox_inst_n461) );
  AOI22X1 aes_core_sbox_inst_U1152 ( .A0(aes_core_sbox_inst_n463), .A1(
        aes_core_sbox_inst_n1720), .B0(aes_core_sbox_inst_n76), .B1(
        aes_core_sbox_inst_n69), .Y(aes_core_sbox_inst_n460) );
  NAND4X1 aes_core_sbox_inst_U1151 ( .A(aes_core_sbox_inst_n411), .B(
        aes_core_sbox_inst_n1706), .C(aes_core_sbox_inst_n460), .D(
        aes_core_sbox_inst_n461), .Y(aes_core_sbox_inst_n441) );
  AOI222X1 aes_core_sbox_inst_U1150 ( .A0(aes_core_sbox_inst_n91), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n101), .B1(
        aes_core_sbox_inst_n96), .C0(aes_core_sbox_inst_n98), .C1(
        aes_core_sbox_inst_n29), .Y(aes_core_sbox_inst_n1056) );
  AOI22X1 aes_core_sbox_inst_U1149 ( .A0(aes_core_sbox_inst_n1058), .A1(
        aes_core_sbox_inst_n24), .B0(aes_core_sbox_inst_n102), .B1(
        aes_core_sbox_inst_n95), .Y(aes_core_sbox_inst_n1055) );
  NAND4X1 aes_core_sbox_inst_U1148 ( .A(aes_core_sbox_inst_n1006), .B(
        aes_core_sbox_inst_n1588), .C(aes_core_sbox_inst_n1055), .D(
        aes_core_sbox_inst_n1056), .Y(aes_core_sbox_inst_n1036) );
  AOI222X1 aes_core_sbox_inst_U1147 ( .A0(aes_core_sbox_inst_n105), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n113), .B1(
        aes_core_sbox_inst_n109), .C0(aes_core_sbox_inst_n630), .C1(
        aes_core_sbox_inst_n19), .Y(aes_core_sbox_inst_n694) );
  AOI22X1 aes_core_sbox_inst_U1146 ( .A0(aes_core_sbox_inst_n696), .A1(
        aes_core_sbox_inst_n243), .B0(aes_core_sbox_inst_n114), .B1(
        aes_core_sbox_inst_n670), .Y(aes_core_sbox_inst_n693) );
  NAND4X1 aes_core_sbox_inst_U1145 ( .A(aes_core_sbox_inst_n644), .B(
        aes_core_sbox_inst_n229), .C(aes_core_sbox_inst_n693), .D(
        aes_core_sbox_inst_n694), .Y(aes_core_sbox_inst_n674) );
  AOI222X1 aes_core_sbox_inst_U1144 ( .A0(aes_core_sbox_inst_n68), .A1(
        aes_core_sbox_inst_n128), .B0(aes_core_sbox_inst_n410), .B1(
        aes_core_sbox_inst_n199), .C0(aes_core_sbox_inst_n74), .C1(
        aes_core_sbox_inst_n140), .Y(aes_core_sbox_inst_n408) );
  NOR2BX1 aes_core_sbox_inst_U1143 ( .AN(aes_core_sbox_inst_n411), .B(
        aes_core_sbox_inst_n76), .Y(aes_core_sbox_inst_n407) );
  NAND4X1 aes_core_sbox_inst_U1142 ( .A(aes_core_sbox_inst_n406), .B(
        aes_core_sbox_inst_n1701), .C(aes_core_sbox_inst_n407), .D(
        aes_core_sbox_inst_n408), .Y(aes_core_sbox_inst_n375) );
  AOI222X1 aes_core_sbox_inst_U1141 ( .A0(aes_core_sbox_inst_n94), .A1(
        aes_core_sbox_inst_n123), .B0(aes_core_sbox_inst_n1005), .B1(
        aes_core_sbox_inst_n174), .C0(aes_core_sbox_inst_n100), .C1(
        aes_core_sbox_inst_n131), .Y(aes_core_sbox_inst_n1003) );
  NOR2BX1 aes_core_sbox_inst_U1140 ( .AN(aes_core_sbox_inst_n1006), .B(
        aes_core_sbox_inst_n102), .Y(aes_core_sbox_inst_n1002) );
  NAND4X1 aes_core_sbox_inst_U1139 ( .A(aes_core_sbox_inst_n1001), .B(
        aes_core_sbox_inst_n1583), .C(aes_core_sbox_inst_n1002), .D(
        aes_core_sbox_inst_n1003), .Y(aes_core_sbox_inst_n970) );
  AOI222X1 aes_core_sbox_inst_U1138 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n3), .B1(
        aes_core_sbox_inst_n69), .C0(aes_core_sbox_inst_n139), .C1(
        aes_core_sbox_inst_n75), .Y(aes_core_sbox_inst_n1165) );
  AOI32X1 aes_core_sbox_inst_U1137 ( .A0(aes_core_sbox_inst_n1732), .A1(
        aes_core_sbox_inst_n49), .A2(aes_core_sbox_inst_n199), .B0(
        aes_core_sbox_inst_n538), .B1(aes_core_sbox_inst_n140), .Y(
        aes_core_sbox_inst_n1164) );
  NAND4X1 aes_core_sbox_inst_U1136 ( .A(aes_core_sbox_inst_n1715), .B(
        aes_core_sbox_inst_n1708), .C(aes_core_sbox_inst_n1164), .D(
        aes_core_sbox_inst_n1165), .Y(aes_core_sbox_inst_n1163) );
  AOI222X1 aes_core_sbox_inst_U1135 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n1045), .B1(
        aes_core_sbox_inst_n95), .C0(aes_core_sbox_inst_n130), .C1(
        aes_core_sbox_inst_n101), .Y(aes_core_sbox_inst_n1269) );
  AOI32X1 aes_core_sbox_inst_U1134 ( .A0(aes_core_sbox_inst_n27), .A1(
        aes_core_sbox_inst_n23), .A2(aes_core_sbox_inst_n174), .B0(
        aes_core_sbox_inst_n1133), .B1(aes_core_sbox_inst_n131), .Y(
        aes_core_sbox_inst_n1268) );
  NAND4X1 aes_core_sbox_inst_U1133 ( .A(aes_core_sbox_inst_n1597), .B(
        aes_core_sbox_inst_n1590), .C(aes_core_sbox_inst_n1268), .D(
        aes_core_sbox_inst_n1269), .Y(aes_core_sbox_inst_n1267) );
  AOI222X1 aes_core_sbox_inst_U1132 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n683), .B1(
        aes_core_sbox_inst_n670), .C0(aes_core_sbox_inst_n135), .C1(
        aes_core_sbox_inst_n113), .Y(aes_core_sbox_inst_n911) );
  AOI32X1 aes_core_sbox_inst_U1131 ( .A0(aes_core_sbox_inst_n18), .A1(
        aes_core_sbox_inst_n15), .A2(aes_core_sbox_inst_n159), .B0(
        aes_core_sbox_inst_n805), .B1(aes_core_sbox_inst_n136), .Y(
        aes_core_sbox_inst_n910) );
  NAND4X1 aes_core_sbox_inst_U1130 ( .A(aes_core_sbox_inst_n238), .B(
        aes_core_sbox_inst_n231), .C(aes_core_sbox_inst_n910), .D(
        aes_core_sbox_inst_n911), .Y(aes_core_sbox_inst_n909) );
  AOI21X1 aes_core_sbox_inst_U1129 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n69), .B0(aes_core_sbox_inst_n477), .Y(
        aes_core_sbox_inst_n1557) );
  AOI222X1 aes_core_sbox_inst_U1128 ( .A0(aes_core_sbox_inst_n68), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n76), .B1(
        aes_core_sbox_inst_n137), .C0(aes_core_sbox_inst_n77), .C1(
        aes_core_sbox_inst_n54), .Y(aes_core_sbox_inst_n1558) );
  NAND4X1 aes_core_sbox_inst_U1127 ( .A(aes_core_sbox_inst_n732), .B(
        aes_core_sbox_inst_n535), .C(aes_core_sbox_inst_n1557), .D(
        aes_core_sbox_inst_n1558), .Y(aes_core_sbox_inst_n1556) );
  AOI21X1 aes_core_sbox_inst_U1126 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n95), .B0(aes_core_sbox_inst_n1072), .Y(
        aes_core_sbox_inst_n1315) );
  AOI222X1 aes_core_sbox_inst_U1125 ( .A0(aes_core_sbox_inst_n94), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n102), .B1(
        aes_core_sbox_inst_n132), .C0(aes_core_sbox_inst_n103), .C1(
        aes_core_sbox_inst_n30), .Y(aes_core_sbox_inst_n1316) );
  NAND4X1 aes_core_sbox_inst_U1124 ( .A(aes_core_sbox_inst_n1237), .B(
        aes_core_sbox_inst_n1130), .C(aes_core_sbox_inst_n1315), .D(
        aes_core_sbox_inst_n1316), .Y(aes_core_sbox_inst_n1314) );
  AOI21X1 aes_core_sbox_inst_U1123 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n670), .B0(aes_core_sbox_inst_n710), .Y(
        aes_core_sbox_inst_n957) );
  AOI222X1 aes_core_sbox_inst_U1122 ( .A0(aes_core_sbox_inst_n108), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n114), .B1(
        aes_core_sbox_inst_n1), .C0(aes_core_sbox_inst_n115), .C1(
        aes_core_sbox_inst_n20), .Y(aes_core_sbox_inst_n958) );
  NAND4X1 aes_core_sbox_inst_U1121 ( .A(aes_core_sbox_inst_n879), .B(
        aes_core_sbox_inst_n802), .C(aes_core_sbox_inst_n957), .D(
        aes_core_sbox_inst_n958), .Y(aes_core_sbox_inst_n956) );
  AOI221X1 aes_core_sbox_inst_U1120 ( .A0(aes_core_sbox_inst_n3), .A1(
        aes_core_sbox_inst_n201), .B0(aes_core_sbox_inst_n469), .B1(
        aes_core_sbox_inst_n139), .C0(aes_core_sbox_inst_n470), .Y(
        aes_core_sbox_inst_n468) );
  AOI222X1 aes_core_sbox_inst_U1119 ( .A0(aes_core_sbox_inst_n471), .A1(
        aes_core_sbox_inst_n49), .B0(aes_core_sbox_inst_n72), .B1(
        aes_core_sbox_inst_n193), .C0(aes_core_sbox_inst_n67), .C1(
        aes_core_sbox_inst_n65), .Y(aes_core_sbox_inst_n467) );
  AOI21X1 aes_core_sbox_inst_U1118 ( .A0(aes_core_sbox_inst_n467), .A1(
        aes_core_sbox_inst_n468), .B0(aes_core_sbox_inst_n1683), .Y(
        aes_core_sbox_inst_n466) );
  AOI221X1 aes_core_sbox_inst_U1117 ( .A0(aes_core_sbox_inst_n1045), .A1(
        aes_core_sbox_inst_n176), .B0(aes_core_sbox_inst_n1064), .B1(
        aes_core_sbox_inst_n130), .C0(aes_core_sbox_inst_n1065), .Y(
        aes_core_sbox_inst_n1063) );
  AOI222X1 aes_core_sbox_inst_U1116 ( .A0(aes_core_sbox_inst_n1066), .A1(
        aes_core_sbox_inst_n23), .B0(aes_core_sbox_inst_n98), .B1(
        aes_core_sbox_inst_n172), .C0(aes_core_sbox_inst_n93), .C1(
        aes_core_sbox_inst_n91), .Y(aes_core_sbox_inst_n1062) );
  AOI21X1 aes_core_sbox_inst_U1115 ( .A0(aes_core_sbox_inst_n1062), .A1(
        aes_core_sbox_inst_n1063), .B0(aes_core_sbox_inst_n617), .Y(
        aes_core_sbox_inst_n1061) );
  AOI221X1 aes_core_sbox_inst_U1114 ( .A0(aes_core_sbox_inst_n683), .A1(
        aes_core_sbox_inst_n162), .B0(aes_core_sbox_inst_n702), .B1(
        aes_core_sbox_inst_n135), .C0(aes_core_sbox_inst_n703), .Y(
        aes_core_sbox_inst_n701) );
  AOI222X1 aes_core_sbox_inst_U1113 ( .A0(aes_core_sbox_inst_n704), .A1(
        aes_core_sbox_inst_n15), .B0(aes_core_sbox_inst_n630), .B1(
        aes_core_sbox_inst_n152), .C0(aes_core_sbox_inst_n107), .C1(
        aes_core_sbox_inst_n105), .Y(aes_core_sbox_inst_n700) );
  AOI21X1 aes_core_sbox_inst_U1112 ( .A0(aes_core_sbox_inst_n700), .A1(
        aes_core_sbox_inst_n701), .B0(aes_core_sbox_inst_n207), .Y(
        aes_core_sbox_inst_n699) );
  AOI22X1 aes_core_sbox_inst_U1111 ( .A0(aes_core_sbox_inst_n742), .A1(
        aes_core_sbox_inst_n127), .B0(aes_core_sbox_inst_n3), .B1(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n1166) );
  AOI222X1 aes_core_sbox_inst_U1110 ( .A0(aes_core_sbox_inst_n69), .A1(
        aes_core_sbox_inst_n75), .B0(aes_core_sbox_inst_n74), .B1(
        aes_core_sbox_inst_n70), .C0(aes_core_sbox_inst_n77), .C1(
        aes_core_sbox_inst_n67), .Y(aes_core_sbox_inst_n1167) );
  NAND4BX1 aes_core_sbox_inst_U1109 ( .AN(aes_core_sbox_inst_n387), .B(
        aes_core_sbox_inst_n1716), .C(aes_core_sbox_inst_n1166), .D(
        aes_core_sbox_inst_n1167), .Y(aes_core_sbox_inst_n1162) );
  AOI22X1 aes_core_sbox_inst_U1108 ( .A0(aes_core_sbox_inst_n1247), .A1(
        aes_core_sbox_inst_n122), .B0(aes_core_sbox_inst_n1045), .B1(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1270) );
  AOI222X1 aes_core_sbox_inst_U1107 ( .A0(aes_core_sbox_inst_n95), .A1(
        aes_core_sbox_inst_n101), .B0(aes_core_sbox_inst_n100), .B1(
        aes_core_sbox_inst_n96), .C0(aes_core_sbox_inst_n103), .C1(
        aes_core_sbox_inst_n93), .Y(aes_core_sbox_inst_n1271) );
  NAND4BX1 aes_core_sbox_inst_U1106 ( .AN(aes_core_sbox_inst_n982), .B(
        aes_core_sbox_inst_n1598), .C(aes_core_sbox_inst_n1270), .D(
        aes_core_sbox_inst_n1271), .Y(aes_core_sbox_inst_n1266) );
  AOI22X1 aes_core_sbox_inst_U1105 ( .A0(aes_core_sbox_inst_n889), .A1(
        aes_core_sbox_inst_n118), .B0(aes_core_sbox_inst_n683), .B1(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n912) );
  AOI222X1 aes_core_sbox_inst_U1104 ( .A0(aes_core_sbox_inst_n670), .A1(
        aes_core_sbox_inst_n113), .B0(aes_core_sbox_inst_n112), .B1(
        aes_core_sbox_inst_n109), .C0(aes_core_sbox_inst_n115), .C1(
        aes_core_sbox_inst_n107), .Y(aes_core_sbox_inst_n913) );
  NAND4BX1 aes_core_sbox_inst_U1103 ( .AN(aes_core_sbox_inst_n620), .B(
        aes_core_sbox_inst_n239), .C(aes_core_sbox_inst_n912), .D(
        aes_core_sbox_inst_n913), .Y(aes_core_sbox_inst_n908) );
  OAI211X1 aes_core_sbox_inst_U1102 ( .A0(aes_core_sbox_inst_n67), .A1(
        aes_core_sbox_inst_n1723), .B0(aes_core_sbox_inst_n600), .C0(
        aes_core_sbox_inst_n601), .Y(aes_core_sbox_inst_n599) );
  AOI222X1 aes_core_sbox_inst_U1101 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n599), .B0(aes_core_sbox_inst_n401), .B1(
        aes_core_sbox_inst_n73), .C0(aes_core_sbox_inst_n573), .C1(
        aes_core_sbox_inst_n192), .Y(aes_core_sbox_inst_n598) );
  AOI21X1 aes_core_sbox_inst_U1100 ( .A0(aes_core_sbox_inst_n603), .A1(
        aes_core_sbox_inst_n6), .B0(aes_core_sbox_inst_n436), .Y(
        aes_core_sbox_inst_n597) );
  NAND4BX1 aes_core_sbox_inst_U1099 ( .AN(aes_core_sbox_inst_n511), .B(
        aes_core_sbox_inst_n581), .C(aes_core_sbox_inst_n597), .D(
        aes_core_sbox_inst_n598), .Y(aes_core_sbox_inst_n566) );
  OAI211X1 aes_core_sbox_inst_U1098 ( .A0(aes_core_sbox_inst_n93), .A1(
        aes_core_sbox_inst_n1605), .B0(aes_core_sbox_inst_n1225), .C0(
        aes_core_sbox_inst_n1226), .Y(aes_core_sbox_inst_n1224) );
  AOI222X1 aes_core_sbox_inst_U1097 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1224), .B0(aes_core_sbox_inst_n996), .B1(
        aes_core_sbox_inst_n99), .C0(aes_core_sbox_inst_n1198), .C1(
        aes_core_sbox_inst_n170), .Y(aes_core_sbox_inst_n1223) );
  AOI21X1 aes_core_sbox_inst_U1096 ( .A0(aes_core_sbox_inst_n1228), .A1(
        aes_core_sbox_inst_n7), .B0(aes_core_sbox_inst_n1031), .Y(
        aes_core_sbox_inst_n1222) );
  NAND4BX1 aes_core_sbox_inst_U1095 ( .AN(aes_core_sbox_inst_n1106), .B(
        aes_core_sbox_inst_n1206), .C(aes_core_sbox_inst_n1222), .D(
        aes_core_sbox_inst_n1223), .Y(aes_core_sbox_inst_n1191) );
  OAI211X1 aes_core_sbox_inst_U1094 ( .A0(aes_core_sbox_inst_n107), .A1(
        aes_core_sbox_inst_n246), .B0(aes_core_sbox_inst_n867), .C0(
        aes_core_sbox_inst_n868), .Y(aes_core_sbox_inst_n866) );
  AOI222X1 aes_core_sbox_inst_U1093 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n866), .B0(aes_core_sbox_inst_n634), .B1(
        aes_core_sbox_inst_n111), .C0(aes_core_sbox_inst_n840), .C1(
        aes_core_sbox_inst_n154), .Y(aes_core_sbox_inst_n865) );
  AOI21X1 aes_core_sbox_inst_U1092 ( .A0(aes_core_sbox_inst_n870), .A1(
        aes_core_sbox_inst_n8), .B0(aes_core_sbox_inst_n669), .Y(
        aes_core_sbox_inst_n864) );
  NAND4BX1 aes_core_sbox_inst_U1091 ( .AN(aes_core_sbox_inst_n778), .B(
        aes_core_sbox_inst_n848), .C(aes_core_sbox_inst_n864), .D(
        aes_core_sbox_inst_n865), .Y(aes_core_sbox_inst_n833) );
  NOR2X1 aes_core_sbox_inst_U1090 ( .A(aes_core_sbox_inst_n15), .B(
        aes_core_sbox_inst_n17), .Y(aes_core_sbox_inst_n635) );
  OAI21X1 aes_core_sbox_inst_U1089 ( .A0(aes_core_sbox_inst_n38), .A1(
        aes_core_sbox_inst_n80), .B0(aes_core_sbox_inst_n144), .Y(
        aes_core_sbox_inst_n1424) );
  AOI21X1 aes_core_sbox_inst_U1088 ( .A0(aes_core_sbox_inst_n293), .A1(
        aes_core_sbox_inst_n1424), .B0(aes_core_sbox_inst_n352), .Y(
        aes_core_sbox_inst_n1417) );
  NAND2X1 aes_core_sbox_inst_U1087 ( .A(aes_core_sbox_inst_n1380), .B(
        aes_core_sbox_inst_n180), .Y(aes_core_sbox_inst_n1429) );
  AOI21X1 aes_core_sbox_inst_U1086 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n489), .Y(
        aes_core_sbox_inst_n744) );
  AOI21X1 aes_core_sbox_inst_U1085 ( .A0(aes_core_sbox_inst_n740), .A1(
        aes_core_sbox_inst_n741), .B0(aes_core_sbox_inst_n1683), .Y(
        aes_core_sbox_inst_n739) );
  NAND4X1 aes_core_sbox_inst_U1084 ( .A(aes_core_sbox_inst_n553), .B(
        aes_core_sbox_inst_n535), .C(aes_core_sbox_inst_n744), .D(
        aes_core_sbox_inst_n745), .Y(aes_core_sbox_inst_n738) );
  AOI21X1 aes_core_sbox_inst_U1083 ( .A0(aes_core_sbox_inst_n529), .A1(
        aes_core_sbox_inst_n738), .B0(aes_core_sbox_inst_n739), .Y(
        aes_core_sbox_inst_n737) );
  AOI21X1 aes_core_sbox_inst_U1082 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n1084), .Y(
        aes_core_sbox_inst_n1249) );
  AOI21X1 aes_core_sbox_inst_U1081 ( .A0(aes_core_sbox_inst_n1245), .A1(
        aes_core_sbox_inst_n1246), .B0(aes_core_sbox_inst_n617), .Y(
        aes_core_sbox_inst_n1244) );
  NAND4X1 aes_core_sbox_inst_U1080 ( .A(aes_core_sbox_inst_n1148), .B(
        aes_core_sbox_inst_n1130), .C(aes_core_sbox_inst_n1249), .D(
        aes_core_sbox_inst_n1250), .Y(aes_core_sbox_inst_n1243) );
  AOI21X1 aes_core_sbox_inst_U1079 ( .A0(aes_core_sbox_inst_n1124), .A1(
        aes_core_sbox_inst_n1243), .B0(aes_core_sbox_inst_n1244), .Y(
        aes_core_sbox_inst_n1242) );
  AOI21X1 aes_core_sbox_inst_U1078 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n722), .Y(
        aes_core_sbox_inst_n891) );
  AOI21X1 aes_core_sbox_inst_U1077 ( .A0(aes_core_sbox_inst_n887), .A1(
        aes_core_sbox_inst_n888), .B0(aes_core_sbox_inst_n207), .Y(
        aes_core_sbox_inst_n886) );
  NAND4X1 aes_core_sbox_inst_U1076 ( .A(aes_core_sbox_inst_n820), .B(
        aes_core_sbox_inst_n802), .C(aes_core_sbox_inst_n891), .D(
        aes_core_sbox_inst_n892), .Y(aes_core_sbox_inst_n885) );
  AOI21X1 aes_core_sbox_inst_U1075 ( .A0(aes_core_sbox_inst_n796), .A1(
        aes_core_sbox_inst_n885), .B0(aes_core_sbox_inst_n886), .Y(
        aes_core_sbox_inst_n884) );
  AOI222X1 aes_core_sbox_inst_U1074 ( .A0(aes_core_sbox_inst_n85), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n272), .B1(
        aes_core_sbox_inst_n43), .C0(aes_core_sbox_inst_n10), .C1(
        aes_core_sbox_inst_n145), .Y(aes_core_sbox_inst_n1527) );
  NAND4X1 aes_core_sbox_inst_U1073 ( .A(aes_core_sbox_inst_n1640), .B(
        aes_core_sbox_inst_n1653), .C(aes_core_sbox_inst_n1348), .D(
        aes_core_sbox_inst_n1529), .Y(aes_core_sbox_inst_n1523) );
  AOI31X1 aes_core_sbox_inst_U1072 ( .A0(aes_core_sbox_inst_n1525), .A1(
        aes_core_sbox_inst_n1526), .A2(aes_core_sbox_inst_n1527), .B0(
        aes_core_sbox_inst_n1624), .Y(aes_core_sbox_inst_n1524) );
  AOI21X1 aes_core_sbox_inst_U1071 ( .A0(aes_core_sbox_inst_n265), .A1(
        aes_core_sbox_inst_n1523), .B0(aes_core_sbox_inst_n1524), .Y(
        aes_core_sbox_inst_n1515) );
  INVX1 aes_core_sbox_inst_U1070 ( .A(aes_core_sbox_inst_n1372), .Y(
        aes_core_sbox_inst_n1625) );
  OAI221X1 aes_core_sbox_inst_U1069 ( .A0(aes_core_sbox_inst_n36), .A1(
        aes_core_sbox_inst_n47), .B0(aes_core_sbox_inst_n45), .B1(
        aes_core_sbox_inst_n32), .C0(aes_core_sbox_inst_n1492), .Y(
        aes_core_sbox_inst_n1487) );
  AOI31X1 aes_core_sbox_inst_U1068 ( .A0(aes_core_sbox_inst_n1489), .A1(
        aes_core_sbox_inst_n1490), .A2(aes_core_sbox_inst_n1491), .B0(
        aes_core_sbox_inst_n1625), .Y(aes_core_sbox_inst_n1488) );
  AOI21X1 aes_core_sbox_inst_U1067 ( .A0(aes_core_sbox_inst_n1374), .A1(
        aes_core_sbox_inst_n1487), .B0(aes_core_sbox_inst_n1488), .Y(
        aes_core_sbox_inst_n1486) );
  AOI31X1 aes_core_sbox_inst_U1066 ( .A0(aes_core_sbox_inst_n383), .A1(
        aes_core_sbox_inst_n49), .A2(aes_core_sbox_inst_n590), .B0(
        aes_core_sbox_inst_n511), .Y(aes_core_sbox_inst_n589) );
  AOI31X1 aes_core_sbox_inst_U1065 ( .A0(aes_core_sbox_inst_n586), .A1(
        aes_core_sbox_inst_n587), .A2(aes_core_sbox_inst_n588), .B0(
        aes_core_sbox_inst_n1687), .Y(aes_core_sbox_inst_n585) );
  OAI221X1 aes_core_sbox_inst_U1064 ( .A0(aes_core_sbox_inst_n202), .A1(
        aes_core_sbox_inst_n1718), .B0(aes_core_sbox_inst_n1709), .B1(
        aes_core_sbox_inst_n128), .C0(aes_core_sbox_inst_n589), .Y(
        aes_core_sbox_inst_n584) );
  AOI21X1 aes_core_sbox_inst_U1063 ( .A0(aes_core_sbox_inst_n440), .A1(
        aes_core_sbox_inst_n584), .B0(aes_core_sbox_inst_n585), .Y(
        aes_core_sbox_inst_n583) );
  AOI31X1 aes_core_sbox_inst_U1062 ( .A0(aes_core_sbox_inst_n978), .A1(
        aes_core_sbox_inst_n23), .A2(aes_core_sbox_inst_n1215), .B0(
        aes_core_sbox_inst_n1106), .Y(aes_core_sbox_inst_n1214) );
  AOI31X1 aes_core_sbox_inst_U1061 ( .A0(aes_core_sbox_inst_n1211), .A1(
        aes_core_sbox_inst_n1212), .A2(aes_core_sbox_inst_n1213), .B0(
        aes_core_sbox_inst_n1569), .Y(aes_core_sbox_inst_n1210) );
  OAI221X1 aes_core_sbox_inst_U1060 ( .A0(aes_core_sbox_inst_n177), .A1(
        aes_core_sbox_inst_n1600), .B0(aes_core_sbox_inst_n1591), .B1(
        aes_core_sbox_inst_n123), .C0(aes_core_sbox_inst_n1214), .Y(
        aes_core_sbox_inst_n1209) );
  AOI21X1 aes_core_sbox_inst_U1059 ( .A0(aes_core_sbox_inst_n1035), .A1(
        aes_core_sbox_inst_n1209), .B0(aes_core_sbox_inst_n1210), .Y(
        aes_core_sbox_inst_n1208) );
  AOI31X1 aes_core_sbox_inst_U1058 ( .A0(aes_core_sbox_inst_n616), .A1(
        aes_core_sbox_inst_n15), .A2(aes_core_sbox_inst_n857), .B0(
        aes_core_sbox_inst_n778), .Y(aes_core_sbox_inst_n856) );
  AOI31X1 aes_core_sbox_inst_U1057 ( .A0(aes_core_sbox_inst_n853), .A1(
        aes_core_sbox_inst_n854), .A2(aes_core_sbox_inst_n855), .B0(
        aes_core_sbox_inst_n211), .Y(aes_core_sbox_inst_n852) );
  OAI221X1 aes_core_sbox_inst_U1056 ( .A0(aes_core_sbox_inst_n163), .A1(
        aes_core_sbox_inst_n16), .B0(aes_core_sbox_inst_n232), .B1(
        aes_core_sbox_inst_n119), .C0(aes_core_sbox_inst_n856), .Y(
        aes_core_sbox_inst_n851) );
  AOI21X1 aes_core_sbox_inst_U1055 ( .A0(aes_core_sbox_inst_n673), .A1(
        aes_core_sbox_inst_n851), .B0(aes_core_sbox_inst_n852), .Y(
        aes_core_sbox_inst_n850) );
  AOI21X1 aes_core_sbox_inst_U1054 ( .A0(aes_core_sbox_inst_n3), .A1(
        aes_core_sbox_inst_n127), .B0(aes_core_sbox_inst_n447), .Y(
        aes_core_sbox_inst_n1549) );
  AOI21X1 aes_core_sbox_inst_U1053 ( .A0(aes_core_sbox_inst_n1045), .A1(
        aes_core_sbox_inst_n122), .B0(aes_core_sbox_inst_n1042), .Y(
        aes_core_sbox_inst_n1307) );
  AOI22X1 aes_core_sbox_inst_U1052 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n127), .B0(aes_core_sbox_inst_n76), .B1(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n600) );
  AOI22X1 aes_core_sbox_inst_U1051 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n122), .B0(aes_core_sbox_inst_n102), .B1(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1225) );
  AOI22X1 aes_core_sbox_inst_U1050 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n118), .B0(aes_core_sbox_inst_n114), .B1(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n867) );
  OAI2BB2X1 aes_core_sbox_inst_U1049 ( .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n1654), .A0N(aes_core_sbox_inst_n45), .A1N(
        aes_core_sbox_inst_n276), .Y(aes_core_sbox_inst_n1454) );
  AOI21X1 aes_core_sbox_inst_U1048 ( .A0(aes_core_sbox_inst_n1718), .A1(
        aes_core_sbox_inst_n1700), .B0(aes_core_sbox_inst_n200), .Y(
        aes_core_sbox_inst_n1179) );
  AOI221X1 aes_core_sbox_inst_U1047 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n67), .B0(aes_core_sbox_inst_n742), .B1(
        aes_core_sbox_inst_n53), .C0(aes_core_sbox_inst_n1179), .Y(
        aes_core_sbox_inst_n1178) );
  AOI222X1 aes_core_sbox_inst_U1046 ( .A0(aes_core_sbox_inst_n139), .A1(
        aes_core_sbox_inst_n73), .B0(aes_core_sbox_inst_n77), .B1(
        aes_core_sbox_inst_n200), .C0(aes_core_sbox_inst_n75), .C1(
        aes_core_sbox_inst_n128), .Y(aes_core_sbox_inst_n1177) );
  AOI21X1 aes_core_sbox_inst_U1045 ( .A0(aes_core_sbox_inst_n1177), .A1(
        aes_core_sbox_inst_n1178), .B0(aes_core_sbox_inst_n1684), .Y(
        aes_core_sbox_inst_n1176) );
  AOI21X1 aes_core_sbox_inst_U1044 ( .A0(aes_core_sbox_inst_n1600), .A1(
        aes_core_sbox_inst_n1582), .B0(aes_core_sbox_inst_n176), .Y(
        aes_core_sbox_inst_n1283) );
  AOI221X1 aes_core_sbox_inst_U1043 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n93), .B0(aes_core_sbox_inst_n1247), .B1(
        aes_core_sbox_inst_n29), .C0(aes_core_sbox_inst_n1283), .Y(
        aes_core_sbox_inst_n1282) );
  AOI222X1 aes_core_sbox_inst_U1042 ( .A0(aes_core_sbox_inst_n130), .A1(
        aes_core_sbox_inst_n99), .B0(aes_core_sbox_inst_n103), .B1(
        aes_core_sbox_inst_n176), .C0(aes_core_sbox_inst_n101), .C1(
        aes_core_sbox_inst_n123), .Y(aes_core_sbox_inst_n1281) );
  AOI21X1 aes_core_sbox_inst_U1041 ( .A0(aes_core_sbox_inst_n1281), .A1(
        aes_core_sbox_inst_n1282), .B0(aes_core_sbox_inst_n1566), .Y(
        aes_core_sbox_inst_n1280) );
  AOI21X1 aes_core_sbox_inst_U1040 ( .A0(aes_core_sbox_inst_n16), .A1(
        aes_core_sbox_inst_n11), .B0(aes_core_sbox_inst_n161), .Y(
        aes_core_sbox_inst_n925) );
  AOI221X1 aes_core_sbox_inst_U1039 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n107), .B0(aes_core_sbox_inst_n889), .B1(
        aes_core_sbox_inst_n19), .C0(aes_core_sbox_inst_n925), .Y(
        aes_core_sbox_inst_n924) );
  AOI222X1 aes_core_sbox_inst_U1038 ( .A0(aes_core_sbox_inst_n135), .A1(
        aes_core_sbox_inst_n111), .B0(aes_core_sbox_inst_n115), .B1(
        aes_core_sbox_inst_n161), .C0(aes_core_sbox_inst_n113), .C1(
        aes_core_sbox_inst_n119), .Y(aes_core_sbox_inst_n923) );
  AOI21X1 aes_core_sbox_inst_U1037 ( .A0(aes_core_sbox_inst_n923), .A1(
        aes_core_sbox_inst_n924), .B0(aes_core_sbox_inst_n208), .Y(
        aes_core_sbox_inst_n922) );
  AOI222X1 aes_core_sbox_inst_U1036 ( .A0(aes_core_sbox_inst_n71), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n3), .B1(
        aes_core_sbox_inst_n194), .C0(aes_core_sbox_inst_n78), .C1(
        aes_core_sbox_inst_n140), .Y(aes_core_sbox_inst_n750) );
  NAND4X1 aes_core_sbox_inst_U1035 ( .A(aes_core_sbox_inst_n1707), .B(
        aes_core_sbox_inst_n553), .C(aes_core_sbox_inst_n411), .D(
        aes_core_sbox_inst_n748), .Y(aes_core_sbox_inst_n747) );
  NAND4BX1 aes_core_sbox_inst_U1034 ( .AN(aes_core_sbox_inst_n448), .B(
        aes_core_sbox_inst_n1707), .C(aes_core_sbox_inst_n749), .D(
        aes_core_sbox_inst_n750), .Y(aes_core_sbox_inst_n746) );
  AOI22X1 aes_core_sbox_inst_U1033 ( .A0(aes_core_sbox_inst_n440), .A1(
        aes_core_sbox_inst_n746), .B0(aes_core_sbox_inst_n592), .B1(
        aes_core_sbox_inst_n747), .Y(aes_core_sbox_inst_n736) );
  AOI222X1 aes_core_sbox_inst_U1032 ( .A0(aes_core_sbox_inst_n97), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n1045), .B1(
        aes_core_sbox_inst_n171), .C0(aes_core_sbox_inst_n104), .C1(
        aes_core_sbox_inst_n131), .Y(aes_core_sbox_inst_n1255) );
  NAND4X1 aes_core_sbox_inst_U1031 ( .A(aes_core_sbox_inst_n1589), .B(
        aes_core_sbox_inst_n1148), .C(aes_core_sbox_inst_n1006), .D(
        aes_core_sbox_inst_n1253), .Y(aes_core_sbox_inst_n1252) );
  NAND4BX1 aes_core_sbox_inst_U1030 ( .AN(aes_core_sbox_inst_n1043), .B(
        aes_core_sbox_inst_n1589), .C(aes_core_sbox_inst_n1254), .D(
        aes_core_sbox_inst_n1255), .Y(aes_core_sbox_inst_n1251) );
  AOI22X1 aes_core_sbox_inst_U1029 ( .A0(aes_core_sbox_inst_n1035), .A1(
        aes_core_sbox_inst_n1251), .B0(aes_core_sbox_inst_n1217), .B1(
        aes_core_sbox_inst_n1252), .Y(aes_core_sbox_inst_n1241) );
  AOI222X1 aes_core_sbox_inst_U1028 ( .A0(aes_core_sbox_inst_n110), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n683), .B1(
        aes_core_sbox_inst_n155), .C0(aes_core_sbox_inst_n116), .C1(
        aes_core_sbox_inst_n136), .Y(aes_core_sbox_inst_n897) );
  NAND4X1 aes_core_sbox_inst_U1027 ( .A(aes_core_sbox_inst_n230), .B(
        aes_core_sbox_inst_n820), .C(aes_core_sbox_inst_n644), .D(
        aes_core_sbox_inst_n895), .Y(aes_core_sbox_inst_n894) );
  NAND4BX1 aes_core_sbox_inst_U1026 ( .AN(aes_core_sbox_inst_n681), .B(
        aes_core_sbox_inst_n230), .C(aes_core_sbox_inst_n896), .D(
        aes_core_sbox_inst_n897), .Y(aes_core_sbox_inst_n893) );
  AOI22X1 aes_core_sbox_inst_U1025 ( .A0(aes_core_sbox_inst_n673), .A1(
        aes_core_sbox_inst_n893), .B0(aes_core_sbox_inst_n859), .B1(
        aes_core_sbox_inst_n894), .Y(aes_core_sbox_inst_n883) );
  AOI222X1 aes_core_sbox_inst_U1024 ( .A0(aes_core_sbox_inst_n383), .A1(
        aes_core_sbox_inst_n1727), .B0(aes_core_sbox_inst_n545), .B1(
        aes_core_sbox_inst_n200), .C0(aes_core_sbox_inst_n76), .C1(
        aes_core_sbox_inst_n54), .Y(aes_core_sbox_inst_n594) );
  NAND4X1 aes_core_sbox_inst_U1023 ( .A(aes_core_sbox_inst_n417), .B(
        aes_core_sbox_inst_n553), .C(aes_core_sbox_inst_n595), .D(
        aes_core_sbox_inst_n596), .Y(aes_core_sbox_inst_n591) );
  NAND4X1 aes_core_sbox_inst_U1022 ( .A(aes_core_sbox_inst_n534), .B(
        aes_core_sbox_inst_n1712), .C(aes_core_sbox_inst_n478), .D(
        aes_core_sbox_inst_n594), .Y(aes_core_sbox_inst_n593) );
  AOI22X1 aes_core_sbox_inst_U1021 ( .A0(aes_core_sbox_inst_n374), .A1(
        aes_core_sbox_inst_n591), .B0(aes_core_sbox_inst_n592), .B1(
        aes_core_sbox_inst_n593), .Y(aes_core_sbox_inst_n582) );
  AOI222X1 aes_core_sbox_inst_U1020 ( .A0(aes_core_sbox_inst_n7), .A1(
        aes_core_sbox_inst_n1609), .B0(aes_core_sbox_inst_n1140), .B1(
        aes_core_sbox_inst_n175), .C0(aes_core_sbox_inst_n102), .C1(
        aes_core_sbox_inst_n30), .Y(aes_core_sbox_inst_n1219) );
  NAND4X1 aes_core_sbox_inst_U1019 ( .A(aes_core_sbox_inst_n1012), .B(
        aes_core_sbox_inst_n1148), .C(aes_core_sbox_inst_n1220), .D(
        aes_core_sbox_inst_n1221), .Y(aes_core_sbox_inst_n1216) );
  NAND4X1 aes_core_sbox_inst_U1018 ( .A(aes_core_sbox_inst_n1129), .B(
        aes_core_sbox_inst_n1594), .C(aes_core_sbox_inst_n1073), .D(
        aes_core_sbox_inst_n1219), .Y(aes_core_sbox_inst_n1218) );
  AOI22X1 aes_core_sbox_inst_U1017 ( .A0(aes_core_sbox_inst_n969), .A1(
        aes_core_sbox_inst_n1216), .B0(aes_core_sbox_inst_n1217), .B1(
        aes_core_sbox_inst_n1218), .Y(aes_core_sbox_inst_n1207) );
  AOI222X1 aes_core_sbox_inst_U1016 ( .A0(aes_core_sbox_inst_n8), .A1(
        aes_core_sbox_inst_n250), .B0(aes_core_sbox_inst_n812), .B1(
        aes_core_sbox_inst_n161), .C0(aes_core_sbox_inst_n114), .C1(
        aes_core_sbox_inst_n20), .Y(aes_core_sbox_inst_n861) );
  NAND4X1 aes_core_sbox_inst_U1015 ( .A(aes_core_sbox_inst_n650), .B(
        aes_core_sbox_inst_n820), .C(aes_core_sbox_inst_n862), .D(
        aes_core_sbox_inst_n863), .Y(aes_core_sbox_inst_n858) );
  NAND4X1 aes_core_sbox_inst_U1014 ( .A(aes_core_sbox_inst_n801), .B(
        aes_core_sbox_inst_n235), .C(aes_core_sbox_inst_n711), .D(
        aes_core_sbox_inst_n861), .Y(aes_core_sbox_inst_n860) );
  AOI22X1 aes_core_sbox_inst_U1013 ( .A0(aes_core_sbox_inst_n607), .A1(
        aes_core_sbox_inst_n858), .B0(aes_core_sbox_inst_n859), .B1(
        aes_core_sbox_inst_n860), .Y(aes_core_sbox_inst_n849) );
  AOI222X1 aes_core_sbox_inst_U1012 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n321), .B0(aes_core_sbox_inst_n90), .B1(
        aes_core_sbox_inst_n43), .C0(aes_core_sbox_inst_n83), .C1(
        aes_core_sbox_inst_n125), .Y(aes_core_sbox_inst_n1520) );
  NAND4X1 aes_core_sbox_inst_U1011 ( .A(aes_core_sbox_inst_n1653), .B(
        aes_core_sbox_inst_n319), .C(aes_core_sbox_inst_n1521), .D(
        aes_core_sbox_inst_n1522), .Y(aes_core_sbox_inst_n1517) );
  OAI211X1 aes_core_sbox_inst_U1010 ( .A0(aes_core_sbox_inst_n1660), .A1(
        aes_core_sbox_inst_n125), .B0(aes_core_sbox_inst_n1519), .C0(
        aes_core_sbox_inst_n1520), .Y(aes_core_sbox_inst_n1518) );
  AOI22X1 aes_core_sbox_inst_U1009 ( .A0(aes_core_sbox_inst_n1372), .A1(
        aes_core_sbox_inst_n1517), .B0(aes_core_sbox_inst_n263), .B1(
        aes_core_sbox_inst_n1518), .Y(aes_core_sbox_inst_n1516) );
  AOI21X1 aes_core_sbox_inst_U1008 ( .A0(aes_core_sbox_inst_n77), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n485), .Y(
        aes_core_sbox_inst_n483) );
  AOI22X1 aes_core_sbox_inst_U1007 ( .A0(aes_core_sbox_inst_n65), .A1(
        aes_core_sbox_inst_n1730), .B0(aes_core_sbox_inst_n54), .B1(
        aes_core_sbox_inst_n50), .Y(aes_core_sbox_inst_n482) );
  OAI22X1 aes_core_sbox_inst_U1006 ( .A0(aes_core_sbox_inst_n186), .A1(
        aes_core_sbox_inst_n482), .B0(aes_core_sbox_inst_n483), .B1(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n481) );
  AOI21X1 aes_core_sbox_inst_U1005 ( .A0(aes_core_sbox_inst_n103), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n1080), .Y(
        aes_core_sbox_inst_n1078) );
  AOI22X1 aes_core_sbox_inst_U1004 ( .A0(aes_core_sbox_inst_n91), .A1(
        aes_core_sbox_inst_n1612), .B0(aes_core_sbox_inst_n1617), .B1(
        aes_core_sbox_inst_n25), .Y(aes_core_sbox_inst_n1077) );
  OAI22X1 aes_core_sbox_inst_U1003 ( .A0(aes_core_sbox_inst_n164), .A1(
        aes_core_sbox_inst_n1077), .B0(aes_core_sbox_inst_n1078), .B1(
        aes_core_sbox_inst_n167), .Y(aes_core_sbox_inst_n1076) );
  AOI22X1 aes_core_sbox_inst_U1002 ( .A0(aes_core_sbox_inst_n105), .A1(
        aes_core_sbox_inst_n253), .B0(aes_core_sbox_inst_n20), .B1(
        aes_core_sbox_inst_n17), .Y(aes_core_sbox_inst_n715) );
  NOR3X1 aes_core_sbox_inst_U1001 ( .A(aes_core_sbox_inst_n49), .B(
        aes_core_sbox_inst_n138), .C(aes_core_sbox_inst_n590), .Y(
        aes_core_sbox_inst_n757) );
  AOI211X1 aes_core_sbox_inst_U1000 ( .A0(aes_core_sbox_inst_n3), .A1(
        aes_core_sbox_inst_n54), .B0(aes_core_sbox_inst_n489), .C0(
        aes_core_sbox_inst_n757), .Y(aes_core_sbox_inst_n756) );
  OAI211X1 aes_core_sbox_inst_U999 ( .A0(aes_core_sbox_inst_n52), .A1(
        aes_core_sbox_inst_n1724), .B0(aes_core_sbox_inst_n432), .C0(
        aes_core_sbox_inst_n756), .Y(aes_core_sbox_inst_n755) );
  AOI22X1 aes_core_sbox_inst_U998 ( .A0(aes_core_sbox_inst_n573), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n186), .B1(
        aes_core_sbox_inst_n755), .Y(aes_core_sbox_inst_n754) );
  NOR3X1 aes_core_sbox_inst_U997 ( .A(aes_core_sbox_inst_n23), .B(
        aes_core_sbox_inst_n129), .C(aes_core_sbox_inst_n1215), .Y(
        aes_core_sbox_inst_n1262) );
  AOI211X1 aes_core_sbox_inst_U996 ( .A0(aes_core_sbox_inst_n1045), .A1(
        aes_core_sbox_inst_n30), .B0(aes_core_sbox_inst_n1084), .C0(
        aes_core_sbox_inst_n1262), .Y(aes_core_sbox_inst_n1261) );
  OAI211X1 aes_core_sbox_inst_U995 ( .A0(aes_core_sbox_inst_n28), .A1(
        aes_core_sbox_inst_n1606), .B0(aes_core_sbox_inst_n1027), .C0(
        aes_core_sbox_inst_n1261), .Y(aes_core_sbox_inst_n1260) );
  AOI22X1 aes_core_sbox_inst_U994 ( .A0(aes_core_sbox_inst_n1198), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n164), .B1(
        aes_core_sbox_inst_n1260), .Y(aes_core_sbox_inst_n1259) );
  NOR3X1 aes_core_sbox_inst_U993 ( .A(aes_core_sbox_inst_n15), .B(
        aes_core_sbox_inst_n134), .C(aes_core_sbox_inst_n857), .Y(
        aes_core_sbox_inst_n904) );
  AOI211X1 aes_core_sbox_inst_U992 ( .A0(aes_core_sbox_inst_n683), .A1(
        aes_core_sbox_inst_n20), .B0(aes_core_sbox_inst_n722), .C0(
        aes_core_sbox_inst_n904), .Y(aes_core_sbox_inst_n903) );
  OAI211X1 aes_core_sbox_inst_U991 ( .A0(aes_core_sbox_inst_n19), .A1(
        aes_core_sbox_inst_n247), .B0(aes_core_sbox_inst_n665), .C0(
        aes_core_sbox_inst_n903), .Y(aes_core_sbox_inst_n902) );
  AOI22X1 aes_core_sbox_inst_U990 ( .A0(aes_core_sbox_inst_n840), .A1(
        aes_core_sbox_inst_n155), .B0(aes_core_sbox_inst_n146), .B1(
        aes_core_sbox_inst_n902), .Y(aes_core_sbox_inst_n901) );
  NOR3X1 aes_core_sbox_inst_U989 ( .A(aes_core_sbox_inst_n34), .B(
        aes_core_sbox_inst_n143), .C(aes_core_sbox_inst_n1334), .Y(
        aes_core_sbox_inst_n1534) );
  AOI211X1 aes_core_sbox_inst_U988 ( .A0(aes_core_sbox_inst_n272), .A1(
        aes_core_sbox_inst_n44), .B0(aes_core_sbox_inst_n1398), .C0(
        aes_core_sbox_inst_n1534), .Y(aes_core_sbox_inst_n1533) );
  AOI21X1 aes_core_sbox_inst_U987 ( .A0(aes_core_sbox_inst_n82), .A1(
        aes_core_sbox_inst_n44), .B0(aes_core_sbox_inst_n1423), .Y(
        aes_core_sbox_inst_n1422) );
  AOI21X1 aes_core_sbox_inst_U986 ( .A0(aes_core_sbox_inst_n1379), .A1(
        aes_core_sbox_inst_n46), .B0(aes_core_sbox_inst_n356), .Y(
        aes_core_sbox_inst_n1421) );
  OAI22X1 aes_core_sbox_inst_U985 ( .A0(aes_core_sbox_inst_n1421), .A1(
        aes_core_sbox_inst_n180), .B0(aes_core_sbox_inst_n179), .B1(
        aes_core_sbox_inst_n1422), .Y(aes_core_sbox_inst_n1419) );
  AOI21X1 aes_core_sbox_inst_U984 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n1735), .B0(aes_core_sbox_inst_n511), .Y(
        aes_core_sbox_inst_n510) );
  AOI21X1 aes_core_sbox_inst_U983 ( .A0(aes_core_sbox_inst_n449), .A1(
        aes_core_sbox_inst_n200), .B0(aes_core_sbox_inst_n68), .Y(
        aes_core_sbox_inst_n509) );
  OAI22X1 aes_core_sbox_inst_U982 ( .A0(aes_core_sbox_inst_n509), .A1(
        aes_core_sbox_inst_n188), .B0(aes_core_sbox_inst_n186), .B1(
        aes_core_sbox_inst_n510), .Y(aes_core_sbox_inst_n505) );
  AOI21X1 aes_core_sbox_inst_U981 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n30), .B0(aes_core_sbox_inst_n1106), .Y(
        aes_core_sbox_inst_n1105) );
  AOI21X1 aes_core_sbox_inst_U980 ( .A0(aes_core_sbox_inst_n1044), .A1(
        aes_core_sbox_inst_n176), .B0(aes_core_sbox_inst_n94), .Y(
        aes_core_sbox_inst_n1104) );
  OAI22X1 aes_core_sbox_inst_U979 ( .A0(aes_core_sbox_inst_n1104), .A1(
        aes_core_sbox_inst_n167), .B0(aes_core_sbox_inst_n164), .B1(
        aes_core_sbox_inst_n1105), .Y(aes_core_sbox_inst_n1100) );
  AOI21X1 aes_core_sbox_inst_U978 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n20), .B0(aes_core_sbox_inst_n778), .Y(
        aes_core_sbox_inst_n777) );
  AOI21X1 aes_core_sbox_inst_U977 ( .A0(aes_core_sbox_inst_n682), .A1(
        aes_core_sbox_inst_n161), .B0(aes_core_sbox_inst_n108), .Y(
        aes_core_sbox_inst_n776) );
  OAI22X1 aes_core_sbox_inst_U976 ( .A0(aes_core_sbox_inst_n776), .A1(
        aes_core_sbox_inst_n148), .B0(aes_core_sbox_inst_n146), .B1(
        aes_core_sbox_inst_n777), .Y(aes_core_sbox_inst_n772) );
  NAND2X1 aes_core_sbox_inst_U975 ( .A(aes_core_sbox_inst_n80), .B(
        aes_core_sbox_inst_n83), .Y(aes_core_sbox_inst_n1339) );
  AOI31X1 aes_core_sbox_inst_U974 ( .A0(aes_core_sbox_inst_n84), .A1(
        aes_core_sbox_inst_n38), .A2(aes_core_sbox_inst_n1357), .B0(
        aes_core_sbox_inst_n1358), .Y(aes_core_sbox_inst_n1349) );
  AOI31X1 aes_core_sbox_inst_U973 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n34), .A2(aes_core_sbox_inst_n1334), .B0(
        aes_core_sbox_inst_n1423), .Y(aes_core_sbox_inst_n1492) );
  INVX1 aes_core_sbox_inst_U972 ( .A(aes_core_sbox_inst_n489), .Y(
        aes_core_sbox_inst_n1722) );
  AOI21X1 aes_core_sbox_inst_U971 ( .A0(aes_core_sbox_inst_n126), .A1(
        aes_core_sbox_inst_n49), .B0(aes_core_sbox_inst_n50), .Y(
        aes_core_sbox_inst_n486) );
  OAI2BB1X1 aes_core_sbox_inst_U970 ( .A0N(aes_core_sbox_inst_n1699), .A1N(
        aes_core_sbox_inst_n1726), .B0(aes_core_sbox_inst_n488), .Y(
        aes_core_sbox_inst_n487) );
  OAI211X1 aes_core_sbox_inst_U969 ( .A0(aes_core_sbox_inst_n486), .A1(
        aes_core_sbox_inst_n1697), .B0(aes_core_sbox_inst_n1722), .C0(
        aes_core_sbox_inst_n487), .Y(aes_core_sbox_inst_n480) );
  AOI21X1 aes_core_sbox_inst_U968 ( .A0(aes_core_sbox_inst_n121), .A1(
        aes_core_sbox_inst_n23), .B0(aes_core_sbox_inst_n25), .Y(
        aes_core_sbox_inst_n1081) );
  OAI2BB1X1 aes_core_sbox_inst_U967 ( .A0N(aes_core_sbox_inst_n1581), .A1N(
        aes_core_sbox_inst_n1608), .B0(aes_core_sbox_inst_n1083), .Y(
        aes_core_sbox_inst_n1082) );
  INVX1 aes_core_sbox_inst_U966 ( .A(aes_core_sbox_inst_n722), .Y(
        aes_core_sbox_inst_n245) );
  AOI21X1 aes_core_sbox_inst_U965 ( .A0(aes_core_sbox_inst_n117), .A1(
        aes_core_sbox_inst_n15), .B0(aes_core_sbox_inst_n17), .Y(
        aes_core_sbox_inst_n719) );
  OAI2BB1X1 aes_core_sbox_inst_U964 ( .A0N(aes_core_sbox_inst_n223), .A1N(
        aes_core_sbox_inst_n249), .B0(aes_core_sbox_inst_n721), .Y(
        aes_core_sbox_inst_n720) );
  OAI211X1 aes_core_sbox_inst_U963 ( .A0(aes_core_sbox_inst_n719), .A1(
        aes_core_sbox_inst_n221), .B0(aes_core_sbox_inst_n245), .C0(
        aes_core_sbox_inst_n720), .Y(aes_core_sbox_inst_n713) );
  AOI211X1 aes_core_sbox_inst_U962 ( .A0(aes_core_sbox_inst_n85), .A1(
        aes_core_sbox_inst_n43), .B0(aes_core_sbox_inst_n1387), .C0(
        aes_core_sbox_inst_n1355), .Y(aes_core_sbox_inst_n1381) );
  OAI2BB1X1 aes_core_sbox_inst_U961 ( .A0N(aes_core_sbox_inst_n1384), .A1N(
        aes_core_sbox_inst_n1385), .B0(aes_core_sbox_inst_n181), .Y(
        aes_core_sbox_inst_n1382) );
  AOI22X1 aes_core_sbox_inst_U960 ( .A0(aes_core_sbox_inst_n291), .A1(
        aes_core_sbox_inst_n84), .B0(aes_core_sbox_inst_n307), .B1(
        aes_core_sbox_inst_n143), .Y(aes_core_sbox_inst_n1383) );
  OAI211X1 aes_core_sbox_inst_U959 ( .A0(aes_core_sbox_inst_n1381), .A1(
        aes_core_sbox_inst_n182), .B0(aes_core_sbox_inst_n1382), .C0(
        aes_core_sbox_inst_n1383), .Y(aes_core_sbox_inst_n1371) );
  AOI222X1 aes_core_sbox_inst_U958 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n90), .B0(aes_core_sbox_inst_n314), .B1(
        aes_core_sbox_inst_n144), .C0(aes_core_sbox_inst_n10), .C1(
        aes_core_sbox_inst_n1677), .Y(aes_core_sbox_inst_n1366) );
  AOI31X1 aes_core_sbox_inst_U957 ( .A0(aes_core_sbox_inst_n1364), .A1(
        aes_core_sbox_inst_n1365), .A2(aes_core_sbox_inst_n1366), .B0(
        aes_core_sbox_inst_n182), .Y(aes_core_sbox_inst_n1360) );
  AOI222X1 aes_core_sbox_inst_U956 ( .A0(aes_core_sbox_inst_n78), .A1(
        aes_core_sbox_inst_n1735), .B0(aes_core_sbox_inst_n410), .B1(
        aes_core_sbox_inst_n140), .C0(aes_core_sbox_inst_n74), .C1(
        aes_core_sbox_inst_n5), .Y(aes_core_sbox_inst_n433) );
  AOI31X1 aes_core_sbox_inst_U955 ( .A0(aes_core_sbox_inst_n431), .A1(
        aes_core_sbox_inst_n432), .A2(aes_core_sbox_inst_n433), .B0(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n427) );
  AOI222X1 aes_core_sbox_inst_U954 ( .A0(aes_core_sbox_inst_n104), .A1(
        aes_core_sbox_inst_n1617), .B0(aes_core_sbox_inst_n1005), .B1(
        aes_core_sbox_inst_n133), .C0(aes_core_sbox_inst_n100), .C1(
        aes_core_sbox_inst_n4), .Y(aes_core_sbox_inst_n1028) );
  AOI31X1 aes_core_sbox_inst_U953 ( .A0(aes_core_sbox_inst_n1026), .A1(
        aes_core_sbox_inst_n1027), .A2(aes_core_sbox_inst_n1028), .B0(
        aes_core_sbox_inst_n166), .Y(aes_core_sbox_inst_n1022) );
  NOR2X1 aes_core_sbox_inst_U952 ( .A(aes_core_sbox_inst_n137), .B(
        aes_core_sbox_inst_n50), .Y(aes_core_sbox_inst_n508) );
  AOI31X1 aes_core_sbox_inst_U951 ( .A0(aes_core_sbox_inst_n502), .A1(
        aes_core_sbox_inst_n535), .A2(aes_core_sbox_inst_n417), .B0(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n1183) );
  AOI31X1 aes_core_sbox_inst_U950 ( .A0(aes_core_sbox_inst_n1187), .A1(
        aes_core_sbox_inst_n476), .A2(aes_core_sbox_inst_n1188), .B0(
        aes_core_sbox_inst_n187), .Y(aes_core_sbox_inst_n1182) );
  AOI21X1 aes_core_sbox_inst_U949 ( .A0(aes_core_sbox_inst_n1185), .A1(
        aes_core_sbox_inst_n1186), .B0(aes_core_sbox_inst_n1691), .Y(
        aes_core_sbox_inst_n1184) );
  OAI31X1 aes_core_sbox_inst_U948 ( .A0(aes_core_sbox_inst_n1182), .A1(
        aes_core_sbox_inst_n1183), .A2(aes_core_sbox_inst_n1184), .B0(
        aes_core_sbox_inst_n1685), .Y(aes_core_sbox_inst_n1173) );
  AOI31X1 aes_core_sbox_inst_U947 ( .A0(aes_core_sbox_inst_n1097), .A1(
        aes_core_sbox_inst_n1130), .A2(aes_core_sbox_inst_n1012), .B0(
        aes_core_sbox_inst_n167), .Y(aes_core_sbox_inst_n1287) );
  AOI31X1 aes_core_sbox_inst_U946 ( .A0(aes_core_sbox_inst_n1291), .A1(
        aes_core_sbox_inst_n1071), .A2(aes_core_sbox_inst_n1292), .B0(
        aes_core_sbox_inst_n165), .Y(aes_core_sbox_inst_n1286) );
  AOI21X1 aes_core_sbox_inst_U945 ( .A0(aes_core_sbox_inst_n1289), .A1(
        aes_core_sbox_inst_n1290), .B0(aes_core_sbox_inst_n1573), .Y(
        aes_core_sbox_inst_n1288) );
  OAI31X1 aes_core_sbox_inst_U944 ( .A0(aes_core_sbox_inst_n1286), .A1(
        aes_core_sbox_inst_n1287), .A2(aes_core_sbox_inst_n1288), .B0(
        aes_core_sbox_inst_n1567), .Y(aes_core_sbox_inst_n1277) );
  NOR2X1 aes_core_sbox_inst_U943 ( .A(aes_core_sbox_inst_n1651), .B(
        aes_core_sbox_inst_n79), .Y(aes_core_sbox_inst_n1356) );
  OAI22X1 aes_core_sbox_inst_U942 ( .A0(aes_core_sbox_inst_n79), .A1(
        aes_core_sbox_inst_n1661), .B0(aes_core_sbox_inst_n44), .B1(
        aes_core_sbox_inst_n1637), .Y(aes_core_sbox_inst_n1387) );
  NAND2X1 aes_core_sbox_inst_U941 ( .A(aes_core_sbox_inst_n293), .B(
        aes_core_sbox_inst_n87), .Y(aes_core_sbox_inst_n338) );
  OAI22X1 aes_core_sbox_inst_U940 ( .A0(aes_core_sbox_inst_n1636), .A1(
        aes_core_sbox_inst_n84), .B0(aes_core_sbox_inst_n31), .B1(
        aes_core_sbox_inst_n1678), .Y(aes_core_sbox_inst_n1367) );
  AOI221X1 aes_core_sbox_inst_U939 ( .A0(aes_core_sbox_inst_n34), .A1(
        aes_core_sbox_inst_n1367), .B0(aes_core_sbox_inst_n356), .B1(
        aes_core_sbox_inst_n1344), .C0(aes_core_sbox_inst_n1368), .Y(
        aes_core_sbox_inst_n1359) );
  AOI222X1 aes_core_sbox_inst_U938 ( .A0(aes_core_sbox_inst_n580), .A1(
        aes_core_sbox_inst_n66), .B0(aes_core_sbox_inst_n77), .B1(
        aes_core_sbox_inst_n139), .C0(aes_core_sbox_inst_n68), .C1(
        aes_core_sbox_inst_n128), .Y(aes_core_sbox_inst_n577) );
  AOI21X1 aes_core_sbox_inst_U937 ( .A0(aes_core_sbox_inst_n1709), .A1(
        aes_core_sbox_inst_n1705), .B0(aes_core_sbox_inst_n187), .Y(
        aes_core_sbox_inst_n575) );
  AOI21X1 aes_core_sbox_inst_U936 ( .A0(aes_core_sbox_inst_n577), .A1(
        aes_core_sbox_inst_n578), .B0(aes_core_sbox_inst_n188), .Y(
        aes_core_sbox_inst_n574) );
  AOI211X1 aes_core_sbox_inst_U935 ( .A0(aes_core_sbox_inst_n573), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n574), .C0(
        aes_core_sbox_inst_n575), .Y(aes_core_sbox_inst_n571) );
  AOI222X1 aes_core_sbox_inst_U934 ( .A0(aes_core_sbox_inst_n1205), .A1(
        aes_core_sbox_inst_n92), .B0(aes_core_sbox_inst_n103), .B1(
        aes_core_sbox_inst_n130), .C0(aes_core_sbox_inst_n94), .C1(
        aes_core_sbox_inst_n123), .Y(aes_core_sbox_inst_n1202) );
  AOI21X1 aes_core_sbox_inst_U933 ( .A0(aes_core_sbox_inst_n1591), .A1(
        aes_core_sbox_inst_n1587), .B0(aes_core_sbox_inst_n165), .Y(
        aes_core_sbox_inst_n1200) );
  AOI21X1 aes_core_sbox_inst_U932 ( .A0(aes_core_sbox_inst_n1202), .A1(
        aes_core_sbox_inst_n1203), .B0(aes_core_sbox_inst_n167), .Y(
        aes_core_sbox_inst_n1199) );
  AOI211X1 aes_core_sbox_inst_U931 ( .A0(aes_core_sbox_inst_n1198), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n1199), .C0(
        aes_core_sbox_inst_n1200), .Y(aes_core_sbox_inst_n1196) );
  AOI222X1 aes_core_sbox_inst_U930 ( .A0(aes_core_sbox_inst_n847), .A1(
        aes_core_sbox_inst_n106), .B0(aes_core_sbox_inst_n115), .B1(
        aes_core_sbox_inst_n135), .C0(aes_core_sbox_inst_n108), .C1(
        aes_core_sbox_inst_n119), .Y(aes_core_sbox_inst_n844) );
  AOI21X1 aes_core_sbox_inst_U929 ( .A0(aes_core_sbox_inst_n232), .A1(
        aes_core_sbox_inst_n228), .B0(aes_core_sbox_inst_n147), .Y(
        aes_core_sbox_inst_n842) );
  AOI21X1 aes_core_sbox_inst_U928 ( .A0(aes_core_sbox_inst_n844), .A1(
        aes_core_sbox_inst_n845), .B0(aes_core_sbox_inst_n148), .Y(
        aes_core_sbox_inst_n841) );
  AOI211X1 aes_core_sbox_inst_U927 ( .A0(aes_core_sbox_inst_n840), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n841), .C0(
        aes_core_sbox_inst_n842), .Y(aes_core_sbox_inst_n838) );
  OAI22X1 aes_core_sbox_inst_U926 ( .A0(aes_core_sbox_inst_n1735), .A1(
        aes_core_sbox_inst_n1723), .B0(aes_core_sbox_inst_n186), .B1(
        aes_core_sbox_inst_n1544), .Y(aes_core_sbox_inst_n1541) );
  OAI221X1 aes_core_sbox_inst_U925 ( .A0(aes_core_sbox_inst_n1703), .A1(
        aes_core_sbox_inst_n53), .B0(aes_core_sbox_inst_n197), .B1(
        aes_core_sbox_inst_n1720), .C0(aes_core_sbox_inst_n518), .Y(
        aes_core_sbox_inst_n1540) );
  OAI32X1 aes_core_sbox_inst_U924 ( .A0(aes_core_sbox_inst_n1732), .A1(
        aes_core_sbox_inst_n1543), .A2(aes_core_sbox_inst_n189), .B0(
        aes_core_sbox_inst_n383), .B1(aes_core_sbox_inst_n1690), .Y(
        aes_core_sbox_inst_n1542) );
  AOI211X1 aes_core_sbox_inst_U923 ( .A0(aes_core_sbox_inst_n404), .A1(
        aes_core_sbox_inst_n1540), .B0(aes_core_sbox_inst_n1541), .C0(
        aes_core_sbox_inst_n1542), .Y(aes_core_sbox_inst_n1539) );
  OAI22X1 aes_core_sbox_inst_U922 ( .A0(aes_core_sbox_inst_n1617), .A1(
        aes_core_sbox_inst_n1605), .B0(aes_core_sbox_inst_n164), .B1(
        aes_core_sbox_inst_n1302), .Y(aes_core_sbox_inst_n1299) );
  OAI221X1 aes_core_sbox_inst_U921 ( .A0(aes_core_sbox_inst_n22), .A1(
        aes_core_sbox_inst_n29), .B0(aes_core_sbox_inst_n174), .B1(
        aes_core_sbox_inst_n24), .C0(aes_core_sbox_inst_n1113), .Y(
        aes_core_sbox_inst_n1298) );
  OAI32X1 aes_core_sbox_inst_U920 ( .A0(aes_core_sbox_inst_n27), .A1(
        aes_core_sbox_inst_n1301), .A2(aes_core_sbox_inst_n167), .B0(
        aes_core_sbox_inst_n978), .B1(aes_core_sbox_inst_n1572), .Y(
        aes_core_sbox_inst_n1300) );
  AOI211X1 aes_core_sbox_inst_U919 ( .A0(aes_core_sbox_inst_n999), .A1(
        aes_core_sbox_inst_n1298), .B0(aes_core_sbox_inst_n1299), .C0(
        aes_core_sbox_inst_n1300), .Y(aes_core_sbox_inst_n1297) );
  OAI22X1 aes_core_sbox_inst_U918 ( .A0(aes_core_sbox_inst_n20), .A1(
        aes_core_sbox_inst_n246), .B0(aes_core_sbox_inst_n146), .B1(
        aes_core_sbox_inst_n944), .Y(aes_core_sbox_inst_n941) );
  OAI221X1 aes_core_sbox_inst_U917 ( .A0(aes_core_sbox_inst_n14), .A1(
        aes_core_sbox_inst_n19), .B0(aes_core_sbox_inst_n160), .B1(
        aes_core_sbox_inst_n243), .C0(aes_core_sbox_inst_n785), .Y(
        aes_core_sbox_inst_n940) );
  OAI32X1 aes_core_sbox_inst_U916 ( .A0(aes_core_sbox_inst_n18), .A1(
        aes_core_sbox_inst_n943), .A2(aes_core_sbox_inst_n148), .B0(
        aes_core_sbox_inst_n8), .B1(aes_core_sbox_inst_n214), .Y(
        aes_core_sbox_inst_n942) );
  AOI211X1 aes_core_sbox_inst_U915 ( .A0(aes_core_sbox_inst_n637), .A1(
        aes_core_sbox_inst_n940), .B0(aes_core_sbox_inst_n941), .C0(
        aes_core_sbox_inst_n942), .Y(aes_core_sbox_inst_n939) );
  AOI21X1 aes_core_sbox_inst_U914 ( .A0(aes_core_sbox_inst_n1656), .A1(
        aes_core_sbox_inst_n40), .B0(aes_core_sbox_inst_n84), .Y(
        aes_core_sbox_inst_n330) );
  OAI22X1 aes_core_sbox_inst_U913 ( .A0(aes_core_sbox_inst_n179), .A1(
        aes_core_sbox_inst_n331), .B0(aes_core_sbox_inst_n332), .B1(
        aes_core_sbox_inst_n31), .Y(aes_core_sbox_inst_n328) );
  OAI32X1 aes_core_sbox_inst_U912 ( .A0(aes_core_sbox_inst_n39), .A1(
        aes_core_sbox_inst_n330), .A2(aes_core_sbox_inst_n181), .B0(
        aes_core_sbox_inst_n80), .B1(aes_core_sbox_inst_n1628), .Y(
        aes_core_sbox_inst_n329) );
  AOI211X1 aes_core_sbox_inst_U911 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n307), .B0(aes_core_sbox_inst_n328), .C0(
        aes_core_sbox_inst_n329), .Y(aes_core_sbox_inst_n326) );
  AOI21X1 aes_core_sbox_inst_U910 ( .A0(aes_core_sbox_inst_n1702), .A1(
        aes_core_sbox_inst_n1723), .B0(aes_core_sbox_inst_n199), .Y(
        aes_core_sbox_inst_n458) );
  AOI31X1 aes_core_sbox_inst_U909 ( .A0(aes_core_sbox_inst_n1732), .A1(
        aes_core_sbox_inst_n49), .A2(aes_core_sbox_inst_n6), .B0(
        aes_core_sbox_inst_n458), .Y(aes_core_sbox_inst_n456) );
  AOI222X1 aes_core_sbox_inst_U908 ( .A0(aes_core_sbox_inst_n65), .A1(
        aes_core_sbox_inst_n1731), .B0(aes_core_sbox_inst_n139), .B1(
        aes_core_sbox_inst_n72), .C0(aes_core_sbox_inst_n69), .C1(
        aes_core_sbox_inst_n73), .Y(aes_core_sbox_inst_n457) );
  OAI211X1 aes_core_sbox_inst_U907 ( .A0(aes_core_sbox_inst_n70), .A1(
        aes_core_sbox_inst_n1700), .B0(aes_core_sbox_inst_n456), .C0(
        aes_core_sbox_inst_n457), .Y(aes_core_sbox_inst_n455) );
  AOI21X1 aes_core_sbox_inst_U906 ( .A0(aes_core_sbox_inst_n1584), .A1(
        aes_core_sbox_inst_n1605), .B0(aes_core_sbox_inst_n174), .Y(
        aes_core_sbox_inst_n1053) );
  AOI31X1 aes_core_sbox_inst_U905 ( .A0(aes_core_sbox_inst_n27), .A1(
        aes_core_sbox_inst_n23), .A2(aes_core_sbox_inst_n978), .B0(
        aes_core_sbox_inst_n1053), .Y(aes_core_sbox_inst_n1051) );
  AOI222X1 aes_core_sbox_inst_U904 ( .A0(aes_core_sbox_inst_n91), .A1(
        aes_core_sbox_inst_n1613), .B0(aes_core_sbox_inst_n130), .B1(
        aes_core_sbox_inst_n98), .C0(aes_core_sbox_inst_n95), .C1(
        aes_core_sbox_inst_n99), .Y(aes_core_sbox_inst_n1052) );
  OAI211X1 aes_core_sbox_inst_U903 ( .A0(aes_core_sbox_inst_n96), .A1(
        aes_core_sbox_inst_n1582), .B0(aes_core_sbox_inst_n1051), .C0(
        aes_core_sbox_inst_n1052), .Y(aes_core_sbox_inst_n1050) );
  AOI21X1 aes_core_sbox_inst_U902 ( .A0(aes_core_sbox_inst_n225), .A1(
        aes_core_sbox_inst_n246), .B0(aes_core_sbox_inst_n159), .Y(
        aes_core_sbox_inst_n691) );
  AOI31X1 aes_core_sbox_inst_U901 ( .A0(aes_core_sbox_inst_n18), .A1(
        aes_core_sbox_inst_n15), .A2(aes_core_sbox_inst_n616), .B0(
        aes_core_sbox_inst_n691), .Y(aes_core_sbox_inst_n689) );
  AOI222X1 aes_core_sbox_inst_U900 ( .A0(aes_core_sbox_inst_n105), .A1(
        aes_core_sbox_inst_n254), .B0(aes_core_sbox_inst_n135), .B1(
        aes_core_sbox_inst_n630), .C0(aes_core_sbox_inst_n670), .C1(
        aes_core_sbox_inst_n111), .Y(aes_core_sbox_inst_n690) );
  OAI211X1 aes_core_sbox_inst_U899 ( .A0(aes_core_sbox_inst_n109), .A1(
        aes_core_sbox_inst_n11), .B0(aes_core_sbox_inst_n689), .C0(
        aes_core_sbox_inst_n690), .Y(aes_core_sbox_inst_n688) );
  OAI221X1 aes_core_sbox_inst_U898 ( .A0(aes_core_sbox_inst_n336), .A1(
        aes_core_sbox_inst_n35), .B0(aes_core_sbox_inst_n37), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n1649), .Y(
        aes_core_sbox_inst_n364) );
  INVX1 aes_core_sbox_inst_U897 ( .A(aes_core_sbox_inst_n10), .Y(
        aes_core_sbox_inst_n1660) );
  INVX1 aes_core_sbox_inst_U896 ( .A(aes_core_sbox_inst_n78), .Y(
        aes_core_sbox_inst_n1723) );
  INVX1 aes_core_sbox_inst_U895 ( .A(aes_core_sbox_inst_n104), .Y(
        aes_core_sbox_inst_n1605) );
  INVX1 aes_core_sbox_inst_U894 ( .A(aes_core_sbox_inst_n116), .Y(
        aes_core_sbox_inst_n246) );
  AOI22X1 aes_core_sbox_inst_U893 ( .A0(aes_core_sbox_inst_n68), .A1(
        aes_core_sbox_inst_n137), .B0(aes_core_sbox_inst_n73), .B1(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n523) );
  OAI2BB1X1 aes_core_sbox_inst_U892 ( .A0N(aes_core_sbox_inst_n66), .A1N(
        aes_core_sbox_inst_n69), .B0(aes_core_sbox_inst_n431), .Y(
        aes_core_sbox_inst_n522) );
  OAI211X1 aes_core_sbox_inst_U891 ( .A0(aes_core_sbox_inst_n1702), .A1(
        aes_core_sbox_inst_n140), .B0(aes_core_sbox_inst_n1717), .C0(
        aes_core_sbox_inst_n523), .Y(aes_core_sbox_inst_n521) );
  AOI222X1 aes_core_sbox_inst_U890 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n521), .B0(aes_core_sbox_inst_n522), .B1(
        aes_core_sbox_inst_n188), .C0(aes_core_sbox_inst_n139), .C1(
        aes_core_sbox_inst_n423), .Y(aes_core_sbox_inst_n520) );
  AOI22X1 aes_core_sbox_inst_U889 ( .A0(aes_core_sbox_inst_n94), .A1(
        aes_core_sbox_inst_n131), .B0(aes_core_sbox_inst_n99), .B1(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n1118) );
  OAI2BB1X1 aes_core_sbox_inst_U888 ( .A0N(aes_core_sbox_inst_n92), .A1N(
        aes_core_sbox_inst_n95), .B0(aes_core_sbox_inst_n1026), .Y(
        aes_core_sbox_inst_n1117) );
  OAI211X1 aes_core_sbox_inst_U887 ( .A0(aes_core_sbox_inst_n1584), .A1(
        aes_core_sbox_inst_n131), .B0(aes_core_sbox_inst_n1599), .C0(
        aes_core_sbox_inst_n1118), .Y(aes_core_sbox_inst_n1116) );
  AOI222X1 aes_core_sbox_inst_U886 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1116), .B0(aes_core_sbox_inst_n1117), .B1(
        aes_core_sbox_inst_n167), .C0(aes_core_sbox_inst_n130), .C1(
        aes_core_sbox_inst_n1018), .Y(aes_core_sbox_inst_n1115) );
  AOI22X1 aes_core_sbox_inst_U885 ( .A0(aes_core_sbox_inst_n108), .A1(
        aes_core_sbox_inst_n136), .B0(aes_core_sbox_inst_n111), .B1(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n790) );
  OAI2BB1X1 aes_core_sbox_inst_U884 ( .A0N(aes_core_sbox_inst_n106), .A1N(
        aes_core_sbox_inst_n670), .B0(aes_core_sbox_inst_n664), .Y(
        aes_core_sbox_inst_n789) );
  OAI211X1 aes_core_sbox_inst_U883 ( .A0(aes_core_sbox_inst_n225), .A1(
        aes_core_sbox_inst_n136), .B0(aes_core_sbox_inst_n240), .C0(
        aes_core_sbox_inst_n790), .Y(aes_core_sbox_inst_n788) );
  AOI222X1 aes_core_sbox_inst_U882 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n788), .B0(aes_core_sbox_inst_n789), .B1(
        aes_core_sbox_inst_n150), .C0(aes_core_sbox_inst_n135), .C1(
        aes_core_sbox_inst_n656), .Y(aes_core_sbox_inst_n787) );
  AOI21X1 aes_core_sbox_inst_U881 ( .A0(aes_core_sbox_inst_n1718), .A1(
        aes_core_sbox_inst_n1706), .B0(aes_core_sbox_inst_n70), .Y(
        aes_core_sbox_inst_n579) );
  AOI211X1 aes_core_sbox_inst_U880 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n192), .B0(aes_core_sbox_inst_n489), .C0(
        aes_core_sbox_inst_n579), .Y(aes_core_sbox_inst_n578) );
  AOI21X1 aes_core_sbox_inst_U879 ( .A0(aes_core_sbox_inst_n1600), .A1(
        aes_core_sbox_inst_n1588), .B0(aes_core_sbox_inst_n96), .Y(
        aes_core_sbox_inst_n1204) );
  AOI211X1 aes_core_sbox_inst_U878 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n170), .B0(aes_core_sbox_inst_n1084), .C0(
        aes_core_sbox_inst_n1204), .Y(aes_core_sbox_inst_n1203) );
  AOI21X1 aes_core_sbox_inst_U877 ( .A0(aes_core_sbox_inst_n16), .A1(
        aes_core_sbox_inst_n229), .B0(aes_core_sbox_inst_n109), .Y(
        aes_core_sbox_inst_n846) );
  AOI211X1 aes_core_sbox_inst_U876 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n154), .B0(aes_core_sbox_inst_n722), .C0(
        aes_core_sbox_inst_n846), .Y(aes_core_sbox_inst_n845) );
  AOI211X1 aes_core_sbox_inst_U875 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n192), .B0(aes_core_sbox_inst_n516), .C0(
        aes_core_sbox_inst_n517), .Y(aes_core_sbox_inst_n514) );
  AOI32X1 aes_core_sbox_inst_U874 ( .A0(aes_core_sbox_inst_n1704), .A1(
        aes_core_sbox_inst_n140), .A2(aes_core_sbox_inst_n399), .B0(
        aes_core_sbox_inst_n1692), .B1(aes_core_sbox_inst_n197), .Y(
        aes_core_sbox_inst_n515) );
  AOI222X1 aes_core_sbox_inst_U873 ( .A0(aes_core_sbox_inst_n65), .A1(
        aes_core_sbox_inst_n1735), .B0(aes_core_sbox_inst_n139), .B1(
        aes_core_sbox_inst_n66), .C0(aes_core_sbox_inst_n67), .C1(
        aes_core_sbox_inst_n71), .Y(aes_core_sbox_inst_n513) );
  OAI221X1 aes_core_sbox_inst_U872 ( .A0(aes_core_sbox_inst_n513), .A1(
        aes_core_sbox_inst_n48), .B0(aes_core_sbox_inst_n514), .B1(
        aes_core_sbox_inst_n190), .C0(aes_core_sbox_inst_n515), .Y(
        aes_core_sbox_inst_n500) );
  AOI211X1 aes_core_sbox_inst_U871 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n170), .B0(aes_core_sbox_inst_n1111), .C0(
        aes_core_sbox_inst_n1112), .Y(aes_core_sbox_inst_n1109) );
  AOI32X1 aes_core_sbox_inst_U870 ( .A0(aes_core_sbox_inst_n1586), .A1(
        aes_core_sbox_inst_n131), .A2(aes_core_sbox_inst_n994), .B0(
        aes_core_sbox_inst_n1574), .B1(aes_core_sbox_inst_n174), .Y(
        aes_core_sbox_inst_n1110) );
  AOI222X1 aes_core_sbox_inst_U869 ( .A0(aes_core_sbox_inst_n91), .A1(
        aes_core_sbox_inst_n1617), .B0(aes_core_sbox_inst_n130), .B1(
        aes_core_sbox_inst_n92), .C0(aes_core_sbox_inst_n93), .C1(
        aes_core_sbox_inst_n97), .Y(aes_core_sbox_inst_n1108) );
  OAI221X1 aes_core_sbox_inst_U868 ( .A0(aes_core_sbox_inst_n1108), .A1(
        aes_core_sbox_inst_n21), .B0(aes_core_sbox_inst_n1109), .B1(
        aes_core_sbox_inst_n166), .C0(aes_core_sbox_inst_n1110), .Y(
        aes_core_sbox_inst_n1095) );
  AOI211X1 aes_core_sbox_inst_U867 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n154), .B0(aes_core_sbox_inst_n783), .C0(
        aes_core_sbox_inst_n784), .Y(aes_core_sbox_inst_n781) );
  AOI32X1 aes_core_sbox_inst_U866 ( .A0(aes_core_sbox_inst_n227), .A1(
        aes_core_sbox_inst_n136), .A2(aes_core_sbox_inst_n632), .B0(
        aes_core_sbox_inst_n216), .B1(aes_core_sbox_inst_n160), .Y(
        aes_core_sbox_inst_n782) );
  AOI222X1 aes_core_sbox_inst_U865 ( .A0(aes_core_sbox_inst_n105), .A1(
        aes_core_sbox_inst_n20), .B0(aes_core_sbox_inst_n135), .B1(
        aes_core_sbox_inst_n106), .C0(aes_core_sbox_inst_n107), .C1(
        aes_core_sbox_inst_n110), .Y(aes_core_sbox_inst_n780) );
  OAI221X1 aes_core_sbox_inst_U864 ( .A0(aes_core_sbox_inst_n780), .A1(
        aes_core_sbox_inst_n13), .B0(aes_core_sbox_inst_n781), .B1(
        aes_core_sbox_inst_n149), .C0(aes_core_sbox_inst_n782), .Y(
        aes_core_sbox_inst_n767) );
  INVX1 aes_core_sbox_inst_U863 ( .A(aes_core_sbox_inst_n1545), .Y(
        aes_core_sbox_inst_n1733) );
  NAND4X1 aes_core_sbox_inst_U862 ( .A(aes_core_sbox_inst_n502), .B(
        aes_core_sbox_inst_n1718), .C(aes_core_sbox_inst_n1564), .D(
        aes_core_sbox_inst_n1565), .Y(aes_core_sbox_inst_n1561) );
  OAI211X1 aes_core_sbox_inst_U861 ( .A0(aes_core_sbox_inst_n1733), .A1(
        aes_core_sbox_inst_n1725), .B0(aes_core_sbox_inst_n419), .C0(
        aes_core_sbox_inst_n416), .Y(aes_core_sbox_inst_n1562) );
  AOI222X1 aes_core_sbox_inst_U860 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n1561), .B0(aes_core_sbox_inst_n1562), .B1(
        aes_core_sbox_inst_n189), .C0(aes_core_sbox_inst_n423), .C1(
        aes_core_sbox_inst_n193), .Y(aes_core_sbox_inst_n1560) );
  INVX1 aes_core_sbox_inst_U859 ( .A(aes_core_sbox_inst_n1303), .Y(
        aes_core_sbox_inst_n1615) );
  NAND4X1 aes_core_sbox_inst_U858 ( .A(aes_core_sbox_inst_n1097), .B(
        aes_core_sbox_inst_n1600), .C(aes_core_sbox_inst_n1322), .D(
        aes_core_sbox_inst_n1323), .Y(aes_core_sbox_inst_n1319) );
  OAI211X1 aes_core_sbox_inst_U857 ( .A0(aes_core_sbox_inst_n1615), .A1(
        aes_core_sbox_inst_n1607), .B0(aes_core_sbox_inst_n1014), .C0(
        aes_core_sbox_inst_n1011), .Y(aes_core_sbox_inst_n1320) );
  AOI222X1 aes_core_sbox_inst_U856 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1319), .B0(aes_core_sbox_inst_n1320), .B1(
        aes_core_sbox_inst_n166), .C0(aes_core_sbox_inst_n1018), .C1(
        aes_core_sbox_inst_n173), .Y(aes_core_sbox_inst_n1318) );
  INVX1 aes_core_sbox_inst_U855 ( .A(aes_core_sbox_inst_n945), .Y(
        aes_core_sbox_inst_n256) );
  NAND4X1 aes_core_sbox_inst_U854 ( .A(aes_core_sbox_inst_n769), .B(
        aes_core_sbox_inst_n16), .C(aes_core_sbox_inst_n964), .D(
        aes_core_sbox_inst_n965), .Y(aes_core_sbox_inst_n961) );
  OAI211X1 aes_core_sbox_inst_U853 ( .A0(aes_core_sbox_inst_n256), .A1(
        aes_core_sbox_inst_n248), .B0(aes_core_sbox_inst_n652), .C0(
        aes_core_sbox_inst_n649), .Y(aes_core_sbox_inst_n962) );
  AOI222X1 aes_core_sbox_inst_U852 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n961), .B0(aes_core_sbox_inst_n962), .B1(
        aes_core_sbox_inst_n148), .C0(aes_core_sbox_inst_n656), .C1(
        aes_core_sbox_inst_n152), .Y(aes_core_sbox_inst_n960) );
  AOI221X1 aes_core_sbox_inst_U851 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n5), .B1(
        aes_core_sbox_inst_n742), .C0(aes_core_sbox_inst_n743), .Y(
        aes_core_sbox_inst_n741) );
  AOI221X1 aes_core_sbox_inst_U850 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n173), .B0(aes_core_sbox_inst_n4), .B1(
        aes_core_sbox_inst_n1247), .C0(aes_core_sbox_inst_n1248), .Y(
        aes_core_sbox_inst_n1246) );
  AOI221X1 aes_core_sbox_inst_U849 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n9), .B1(
        aes_core_sbox_inst_n889), .C0(aes_core_sbox_inst_n890), .Y(
        aes_core_sbox_inst_n888) );
  AOI211X1 aes_core_sbox_inst_U848 ( .A0(aes_core_sbox_inst_n75), .A1(
        aes_core_sbox_inst_n128), .B0(aes_core_sbox_inst_n421), .C0(
        aes_core_sbox_inst_n563), .Y(aes_core_sbox_inst_n556) );
  NOR4BX1 aes_core_sbox_inst_U847 ( .AN(aes_core_sbox_inst_n559), .B(
        aes_core_sbox_inst_n447), .C(aes_core_sbox_inst_n560), .D(
        aes_core_sbox_inst_n469), .Y(aes_core_sbox_inst_n558) );
  AOI211X1 aes_core_sbox_inst_U846 ( .A0(aes_core_sbox_inst_n139), .A1(
        aes_core_sbox_inst_n49), .B0(aes_core_sbox_inst_n562), .C0(
        aes_core_sbox_inst_n73), .Y(aes_core_sbox_inst_n557) );
  OAI222X1 aes_core_sbox_inst_U845 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n556), .B0(aes_core_sbox_inst_n557), .B1(
        aes_core_sbox_inst_n48), .C0(aes_core_sbox_inst_n558), .C1(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n547) );
  AOI211X1 aes_core_sbox_inst_U844 ( .A0(aes_core_sbox_inst_n101), .A1(
        aes_core_sbox_inst_n123), .B0(aes_core_sbox_inst_n1016), .C0(
        aes_core_sbox_inst_n1158), .Y(aes_core_sbox_inst_n1151) );
  NOR4BX1 aes_core_sbox_inst_U843 ( .AN(aes_core_sbox_inst_n1154), .B(
        aes_core_sbox_inst_n1042), .C(aes_core_sbox_inst_n1155), .D(
        aes_core_sbox_inst_n1064), .Y(aes_core_sbox_inst_n1153) );
  AOI211X1 aes_core_sbox_inst_U842 ( .A0(aes_core_sbox_inst_n130), .A1(
        aes_core_sbox_inst_n23), .B0(aes_core_sbox_inst_n1157), .C0(
        aes_core_sbox_inst_n99), .Y(aes_core_sbox_inst_n1152) );
  OAI222X1 aes_core_sbox_inst_U841 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1151), .B0(aes_core_sbox_inst_n1152), .B1(
        aes_core_sbox_inst_n21), .C0(aes_core_sbox_inst_n1153), .C1(
        aes_core_sbox_inst_n166), .Y(aes_core_sbox_inst_n1142) );
  AOI211X1 aes_core_sbox_inst_U840 ( .A0(aes_core_sbox_inst_n113), .A1(
        aes_core_sbox_inst_n119), .B0(aes_core_sbox_inst_n654), .C0(
        aes_core_sbox_inst_n830), .Y(aes_core_sbox_inst_n823) );
  NOR4BX1 aes_core_sbox_inst_U839 ( .AN(aes_core_sbox_inst_n826), .B(
        aes_core_sbox_inst_n680), .C(aes_core_sbox_inst_n827), .D(
        aes_core_sbox_inst_n702), .Y(aes_core_sbox_inst_n825) );
  AOI211X1 aes_core_sbox_inst_U838 ( .A0(aes_core_sbox_inst_n135), .A1(
        aes_core_sbox_inst_n15), .B0(aes_core_sbox_inst_n829), .C0(
        aes_core_sbox_inst_n111), .Y(aes_core_sbox_inst_n824) );
  OAI222X1 aes_core_sbox_inst_U837 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n823), .B0(aes_core_sbox_inst_n824), .B1(
        aes_core_sbox_inst_n13), .C0(aes_core_sbox_inst_n825), .C1(
        aes_core_sbox_inst_n150), .Y(aes_core_sbox_inst_n814) );
  INVX1 aes_core_sbox_inst_U836 ( .A(aes_core_sbox_inst_n318), .Y(
        aes_core_sbox_inst_n1643) );
  AOI221X1 aes_core_sbox_inst_U835 ( .A0(aes_core_sbox_inst_n321), .A1(
        aes_core_sbox_inst_n47), .B0(aes_core_sbox_inst_n82), .B1(
        aes_core_sbox_inst_n41), .C0(aes_core_sbox_inst_n322), .Y(
        aes_core_sbox_inst_n308) );
  OAI222X1 aes_core_sbox_inst_U834 ( .A0(aes_core_sbox_inst_n308), .A1(
        aes_core_sbox_inst_n1630), .B0(aes_core_sbox_inst_n1643), .B1(
        aes_core_sbox_inst_n181), .C0(aes_core_sbox_inst_n179), .C1(
        aes_core_sbox_inst_n309), .Y(aes_core_sbox_inst_n297) );
  INVX1 aes_core_sbox_inst_U833 ( .A(aes_core_sbox_inst_n735), .Y(
        aes_core_sbox_inst_n1719) );
  AOI221X1 aes_core_sbox_inst_U832 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n68), .B1(
        aes_core_sbox_inst_n194), .C0(aes_core_sbox_inst_n1719), .Y(
        aes_core_sbox_inst_n745) );
  AOI21X1 aes_core_sbox_inst_U831 ( .A0(aes_core_sbox_inst_n1720), .A1(
        aes_core_sbox_inst_n1698), .B0(aes_core_sbox_inst_n193), .Y(
        aes_core_sbox_inst_n734) );
  AOI221X1 aes_core_sbox_inst_U830 ( .A0(aes_core_sbox_inst_n74), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n545), .B1(
        aes_core_sbox_inst_n6), .C0(aes_core_sbox_inst_n734), .Y(
        aes_core_sbox_inst_n733) );
  INVX1 aes_core_sbox_inst_U829 ( .A(aes_core_sbox_inst_n1240), .Y(
        aes_core_sbox_inst_n1601) );
  AOI221X1 aes_core_sbox_inst_U828 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n94), .B1(
        aes_core_sbox_inst_n171), .C0(aes_core_sbox_inst_n1601), .Y(
        aes_core_sbox_inst_n1250) );
  AOI21X1 aes_core_sbox_inst_U827 ( .A0(aes_core_sbox_inst_n24), .A1(
        aes_core_sbox_inst_n1580), .B0(aes_core_sbox_inst_n171), .Y(
        aes_core_sbox_inst_n1239) );
  AOI221X1 aes_core_sbox_inst_U826 ( .A0(aes_core_sbox_inst_n100), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n1140), .B1(
        aes_core_sbox_inst_n7), .C0(aes_core_sbox_inst_n1239), .Y(
        aes_core_sbox_inst_n1238) );
  INVX1 aes_core_sbox_inst_U825 ( .A(aes_core_sbox_inst_n882), .Y(
        aes_core_sbox_inst_n242) );
  AOI221X1 aes_core_sbox_inst_U824 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n108), .B1(
        aes_core_sbox_inst_n152), .C0(aes_core_sbox_inst_n242), .Y(
        aes_core_sbox_inst_n892) );
  AOI21X1 aes_core_sbox_inst_U823 ( .A0(aes_core_sbox_inst_n243), .A1(
        aes_core_sbox_inst_n222), .B0(aes_core_sbox_inst_n153), .Y(
        aes_core_sbox_inst_n881) );
  AOI221X1 aes_core_sbox_inst_U822 ( .A0(aes_core_sbox_inst_n112), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n812), .B1(
        aes_core_sbox_inst_n8), .C0(aes_core_sbox_inst_n881), .Y(
        aes_core_sbox_inst_n880) );
  AOI211X1 aes_core_sbox_inst_U821 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n194), .B0(aes_core_sbox_inst_n542), .C0(
        aes_core_sbox_inst_n543), .Y(aes_core_sbox_inst_n541) );
  AOI211X1 aes_core_sbox_inst_U820 ( .A0(aes_core_sbox_inst_n545), .A1(
        aes_core_sbox_inst_n199), .B0(aes_core_sbox_inst_n546), .C0(
        aes_core_sbox_inst_n68), .Y(aes_core_sbox_inst_n539) );
  AOI21X1 aes_core_sbox_inst_U819 ( .A0(aes_core_sbox_inst_n71), .A1(
        aes_core_sbox_inst_n127), .B0(aes_core_sbox_inst_n430), .Y(
        aes_core_sbox_inst_n540) );
  OAI222X1 aes_core_sbox_inst_U818 ( .A0(aes_core_sbox_inst_n539), .A1(
        aes_core_sbox_inst_n188), .B0(aes_core_sbox_inst_n540), .B1(
        aes_core_sbox_inst_n1691), .C0(aes_core_sbox_inst_n187), .C1(
        aes_core_sbox_inst_n541), .Y(aes_core_sbox_inst_n528) );
  AOI211X1 aes_core_sbox_inst_U817 ( .A0(aes_core_sbox_inst_n102), .A1(
        aes_core_sbox_inst_n172), .B0(aes_core_sbox_inst_n1137), .C0(
        aes_core_sbox_inst_n1138), .Y(aes_core_sbox_inst_n1136) );
  AOI211X1 aes_core_sbox_inst_U816 ( .A0(aes_core_sbox_inst_n1140), .A1(
        aes_core_sbox_inst_n174), .B0(aes_core_sbox_inst_n1141), .C0(
        aes_core_sbox_inst_n94), .Y(aes_core_sbox_inst_n1134) );
  AOI21X1 aes_core_sbox_inst_U815 ( .A0(aes_core_sbox_inst_n97), .A1(
        aes_core_sbox_inst_n122), .B0(aes_core_sbox_inst_n1025), .Y(
        aes_core_sbox_inst_n1135) );
  OAI222X1 aes_core_sbox_inst_U814 ( .A0(aes_core_sbox_inst_n1134), .A1(
        aes_core_sbox_inst_n167), .B0(aes_core_sbox_inst_n1135), .B1(
        aes_core_sbox_inst_n1573), .C0(aes_core_sbox_inst_n165), .C1(
        aes_core_sbox_inst_n1136), .Y(aes_core_sbox_inst_n1123) );
  AOI211X1 aes_core_sbox_inst_U813 ( .A0(aes_core_sbox_inst_n114), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n809), .C0(
        aes_core_sbox_inst_n810), .Y(aes_core_sbox_inst_n808) );
  AOI211X1 aes_core_sbox_inst_U812 ( .A0(aes_core_sbox_inst_n812), .A1(
        aes_core_sbox_inst_n160), .B0(aes_core_sbox_inst_n813), .C0(
        aes_core_sbox_inst_n108), .Y(aes_core_sbox_inst_n806) );
  AOI21X1 aes_core_sbox_inst_U811 ( .A0(aes_core_sbox_inst_n110), .A1(
        aes_core_sbox_inst_n118), .B0(aes_core_sbox_inst_n663), .Y(
        aes_core_sbox_inst_n807) );
  OAI222X1 aes_core_sbox_inst_U810 ( .A0(aes_core_sbox_inst_n806), .A1(
        aes_core_sbox_inst_n148), .B0(aes_core_sbox_inst_n807), .B1(
        aes_core_sbox_inst_n215), .C0(aes_core_sbox_inst_n147), .C1(
        aes_core_sbox_inst_n808), .Y(aes_core_sbox_inst_n795) );
  AOI222X1 aes_core_sbox_inst_U809 ( .A0(aes_core_sbox_inst_n139), .A1(
        aes_core_sbox_inst_n66), .B0(aes_core_sbox_inst_n78), .B1(
        aes_core_sbox_inst_n53), .C0(aes_core_sbox_inst_n77), .C1(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n740) );
  AOI222X1 aes_core_sbox_inst_U808 ( .A0(aes_core_sbox_inst_n130), .A1(
        aes_core_sbox_inst_n92), .B0(aes_core_sbox_inst_n104), .B1(
        aes_core_sbox_inst_n29), .C0(aes_core_sbox_inst_n103), .C1(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1245) );
  AOI222X1 aes_core_sbox_inst_U807 ( .A0(aes_core_sbox_inst_n135), .A1(
        aes_core_sbox_inst_n106), .B0(aes_core_sbox_inst_n116), .B1(
        aes_core_sbox_inst_n19), .C0(aes_core_sbox_inst_n115), .C1(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n887) );
  INVX1 aes_core_sbox_inst_U806 ( .A(aes_core_sbox_inst_n1364), .Y(
        aes_core_sbox_inst_n1652) );
  AOI211X1 aes_core_sbox_inst_U805 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n88), .B0(aes_core_sbox_inst_n1437), .C0(
        aes_core_sbox_inst_n1432), .Y(aes_core_sbox_inst_n1436) );
  AOI21X1 aes_core_sbox_inst_U804 ( .A0(aes_core_sbox_inst_n84), .A1(
        aes_core_sbox_inst_n321), .B0(aes_core_sbox_inst_n1652), .Y(
        aes_core_sbox_inst_n1435) );
  OAI222X1 aes_core_sbox_inst_U803 ( .A0(aes_core_sbox_inst_n2), .A1(
        aes_core_sbox_inst_n1632), .B0(aes_core_sbox_inst_n179), .B1(
        aes_core_sbox_inst_n1435), .C0(aes_core_sbox_inst_n1436), .C1(
        aes_core_sbox_inst_n181), .Y(aes_core_sbox_inst_n1434) );
  AOI211X1 aes_core_sbox_inst_U802 ( .A0(aes_core_sbox_inst_n111), .A1(
        aes_core_sbox_inst_n136), .B0(aes_core_sbox_inst_n654), .C0(
        aes_core_sbox_inst_n655), .Y(aes_core_sbox_inst_n651) );
  INVX1 aes_core_sbox_inst_U801 ( .A(aes_core_sbox_inst_n656), .Y(
        aes_core_sbox_inst_n217) );
  OAI222X1 aes_core_sbox_inst_U800 ( .A0(aes_core_sbox_inst_n109), .A1(
        aes_core_sbox_inst_n217), .B0(aes_core_sbox_inst_n651), .B1(
        aes_core_sbox_inst_n149), .C0(aes_core_sbox_inst_n215), .C1(
        aes_core_sbox_inst_n652), .Y(aes_core_sbox_inst_n646) );
  AOI211X1 aes_core_sbox_inst_U799 ( .A0(aes_core_sbox_inst_n80), .A1(
        aes_core_sbox_inst_n86), .B0(aes_core_sbox_inst_n1355), .C0(
        aes_core_sbox_inst_n267), .Y(aes_core_sbox_inst_n1354) );
  AOI221X1 aes_core_sbox_inst_U798 ( .A0(aes_core_sbox_inst_n79), .A1(
        aes_core_sbox_inst_n87), .B0(aes_core_sbox_inst_n82), .B1(
        aes_core_sbox_inst_n145), .C0(aes_core_sbox_inst_n1356), .Y(
        aes_core_sbox_inst_n1353) );
  OAI222X1 aes_core_sbox_inst_U797 ( .A0(aes_core_sbox_inst_n1353), .A1(
        aes_core_sbox_inst_n181), .B0(aes_core_sbox_inst_n184), .B1(
        aes_core_sbox_inst_n1354), .C0(aes_core_sbox_inst_n125), .C1(
        aes_core_sbox_inst_n1632), .Y(aes_core_sbox_inst_n1350) );
  INVX1 aes_core_sbox_inst_U796 ( .A(aes_core_sbox_inst_n272), .Y(
        aes_core_sbox_inst_n1654) );
  AOI222X1 aes_core_sbox_inst_U795 ( .A0(aes_core_sbox_inst_n65), .A1(
        aes_core_sbox_inst_n1731), .B0(aes_core_sbox_inst_n78), .B1(
        aes_core_sbox_inst_n199), .C0(aes_core_sbox_inst_n75), .C1(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n596) );
  AOI222X1 aes_core_sbox_inst_U794 ( .A0(aes_core_sbox_inst_n91), .A1(
        aes_core_sbox_inst_n1613), .B0(aes_core_sbox_inst_n104), .B1(
        aes_core_sbox_inst_n174), .C0(aes_core_sbox_inst_n101), .C1(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1221) );
  AOI222X1 aes_core_sbox_inst_U793 ( .A0(aes_core_sbox_inst_n105), .A1(
        aes_core_sbox_inst_n254), .B0(aes_core_sbox_inst_n116), .B1(
        aes_core_sbox_inst_n159), .C0(aes_core_sbox_inst_n113), .C1(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n863) );
  INVX1 aes_core_sbox_inst_U792 ( .A(aes_core_sbox_inst_n1357), .Y(
        aes_core_sbox_inst_n1630) );
  NOR2X1 aes_core_sbox_inst_U791 ( .A(aes_core_sbox_inst_n49), .B(
        aes_core_sbox_inst_n50), .Y(aes_core_sbox_inst_n402) );
  NOR2X1 aes_core_sbox_inst_U790 ( .A(aes_core_sbox_inst_n23), .B(
        aes_core_sbox_inst_n25), .Y(aes_core_sbox_inst_n997) );
  BUFX3 aes_core_sbox_inst_U789 ( .A(aes_core_sbox_inst_n997), .Y(
        aes_core_sbox_inst_n91) );
  AOI211X1 aes_core_sbox_inst_U788 ( .A0(aes_core_sbox_inst_n73), .A1(
        aes_core_sbox_inst_n140), .B0(aes_core_sbox_inst_n421), .C0(
        aes_core_sbox_inst_n422), .Y(aes_core_sbox_inst_n418) );
  INVX1 aes_core_sbox_inst_U787 ( .A(aes_core_sbox_inst_n423), .Y(
        aes_core_sbox_inst_n1693) );
  OAI222X1 aes_core_sbox_inst_U786 ( .A0(aes_core_sbox_inst_n70), .A1(
        aes_core_sbox_inst_n1693), .B0(aes_core_sbox_inst_n418), .B1(
        aes_core_sbox_inst_n188), .C0(aes_core_sbox_inst_n1691), .C1(
        aes_core_sbox_inst_n419), .Y(aes_core_sbox_inst_n413) );
  AOI211X1 aes_core_sbox_inst_U785 ( .A0(aes_core_sbox_inst_n99), .A1(
        aes_core_sbox_inst_n131), .B0(aes_core_sbox_inst_n1016), .C0(
        aes_core_sbox_inst_n1017), .Y(aes_core_sbox_inst_n1013) );
  INVX1 aes_core_sbox_inst_U784 ( .A(aes_core_sbox_inst_n1018), .Y(
        aes_core_sbox_inst_n1575) );
  OAI222X1 aes_core_sbox_inst_U783 ( .A0(aes_core_sbox_inst_n96), .A1(
        aes_core_sbox_inst_n1575), .B0(aes_core_sbox_inst_n1013), .B1(
        aes_core_sbox_inst_n167), .C0(aes_core_sbox_inst_n1573), .C1(
        aes_core_sbox_inst_n1014), .Y(aes_core_sbox_inst_n1008) );
  INVX1 aes_core_sbox_inst_U782 ( .A(aes_core_sbox_inst_n186), .Y(
        aes_core_sbox_inst_n188) );
  INVX1 aes_core_sbox_inst_U781 ( .A(aes_core_sbox_inst_n159), .Y(
        aes_core_sbox_inst_n161) );
  INVX1 aes_core_sbox_inst_U780 ( .A(aes_core_n3), .Y(aes_core_sbox_inst_n194)
         );
  INVX1 aes_core_sbox_inst_U779 ( .A(aes_core_sbox_inst_n164), .Y(
        aes_core_sbox_inst_n167) );
  INVX1 aes_core_sbox_inst_U778 ( .A(aes_core_sbox_inst_n184), .Y(
        aes_core_sbox_inst_n181) );
  INVX1 aes_core_sbox_inst_U777 ( .A(aes_core_sbox_inst_n164), .Y(
        aes_core_sbox_inst_n166) );
  INVX1 aes_core_sbox_inst_U776 ( .A(aes_core_sbox_inst_n154), .Y(
        aes_core_sbox_inst_n152) );
  INVX1 aes_core_sbox_inst_U775 ( .A(aes_core_sbox_inst_n199), .Y(
        aes_core_sbox_inst_n200) );
  INVX1 aes_core_sbox_inst_U774 ( .A(aes_core_sbox_inst_n192), .Y(
        aes_core_sbox_inst_n193) );
  INVX1 aes_core_sbox_inst_U773 ( .A(aes_core_sbox_inst_n184), .Y(
        aes_core_sbox_inst_n180) );
  INVX1 aes_core_sbox_inst_U772 ( .A(aes_core_sbox_inst_n146), .Y(
        aes_core_sbox_inst_n148) );
  INVX1 aes_core_sbox_inst_U771 ( .A(aes_core_sbox_inst_n163), .Y(
        aes_core_sbox_inst_n160) );
  BUFX3 aes_core_sbox_inst_U770 ( .A(aes_core_sbox_inst_n1678), .Y(
        aes_core_sbox_inst_n45) );
  INVX1 aes_core_sbox_inst_U769 ( .A(aes_core_sbox_inst_n1471), .Y(
        aes_core_sbox_inst_n1618) );
  INVX1 aes_core_sbox_inst_U768 ( .A(aes_core_sbox_inst_n374), .Y(
        aes_core_sbox_inst_n1683) );
  INVX1 aes_core_sbox_inst_U767 ( .A(aes_core_sbox_inst_n969), .Y(
        aes_core_sbox_inst_n617) );
  INVX1 aes_core_sbox_inst_U766 ( .A(aes_core_sbox_inst_n607), .Y(
        aes_core_sbox_inst_n207) );
  NOR2X1 aes_core_sbox_inst_U765 ( .A(aes_core_sbox_inst_n18), .B(
        aes_core_sbox_inst_n15), .Y(aes_core_sbox_inst_n702) );
  INVX1 aes_core_sbox_inst_U764 ( .A(aes_core_sbox_inst_n751), .Y(
        aes_core_sbox_inst_n1692) );
  INVX1 aes_core_sbox_inst_U763 ( .A(aes_core_sbox_inst_n1256), .Y(
        aes_core_sbox_inst_n1574) );
  INVX1 aes_core_sbox_inst_U762 ( .A(aes_core_sbox_inst_n898), .Y(
        aes_core_sbox_inst_n216) );
  INVX1 aes_core_sbox_inst_U761 ( .A(aes_core_sbox_inst_n775), .Y(
        aes_core_sbox_inst_n249) );
  AOI2BB1X1 aes_core_sbox_inst_U760 ( .A0N(aes_core_sbox_inst_n87), .A1N(
        aes_core_sbox_inst_n1379), .B0(aes_core_sbox_inst_n143), .Y(
        aes_core_sbox_inst_n1469) );
  AOI2BB1X1 aes_core_sbox_inst_U759 ( .A0N(aes_core_sbox_inst_n65), .A1N(
        aes_core_sbox_inst_n449), .B0(aes_core_sbox_inst_n138), .Y(
        aes_core_sbox_inst_n560) );
  AOI2BB1X1 aes_core_sbox_inst_U758 ( .A0N(aes_core_sbox_inst_n91), .A1N(
        aes_core_sbox_inst_n1044), .B0(aes_core_sbox_inst_n129), .Y(
        aes_core_sbox_inst_n1155) );
  AOI2BB1X1 aes_core_sbox_inst_U757 ( .A0N(aes_core_sbox_inst_n105), .A1N(
        aes_core_sbox_inst_n682), .B0(aes_core_sbox_inst_n134), .Y(
        aes_core_sbox_inst_n827) );
  NAND3X1 aes_core_sbox_inst_U756 ( .A(aes_core_sbox_inst_n127), .B(
        aes_core_sbox_inst_n49), .C(aes_core_sbox_inst_n590), .Y(
        aes_core_sbox_inst_n595) );
  NAND3X1 aes_core_sbox_inst_U755 ( .A(aes_core_sbox_inst_n122), .B(
        aes_core_sbox_inst_n23), .C(aes_core_sbox_inst_n1215), .Y(
        aes_core_sbox_inst_n1220) );
  NAND3X1 aes_core_sbox_inst_U754 ( .A(aes_core_sbox_inst_n118), .B(
        aes_core_sbox_inst_n15), .C(aes_core_sbox_inst_n857), .Y(
        aes_core_sbox_inst_n862) );
  INVX1 aes_core_sbox_inst_U753 ( .A(aes_core_sbox_inst_n590), .Y(
        aes_core_sbox_inst_n1727) );
  INVX1 aes_core_sbox_inst_U752 ( .A(aes_core_sbox_inst_n1215), .Y(
        aes_core_sbox_inst_n1609) );
  INVX1 aes_core_sbox_inst_U751 ( .A(aes_core_sbox_inst_n857), .Y(
        aes_core_sbox_inst_n250) );
  OAI22X1 aes_core_sbox_inst_U750 ( .A0(aes_core_sbox_inst_n143), .A1(
        aes_core_sbox_inst_n32), .B0(aes_core_sbox_inst_n46), .B1(
        aes_core_sbox_inst_n1651), .Y(aes_core_sbox_inst_n289) );
  AOI22X1 aes_core_sbox_inst_U749 ( .A0(aes_core_sbox_inst_n179), .A1(
        aes_core_sbox_inst_n289), .B0(aes_core_sbox_inst_n290), .B1(
        aes_core_sbox_inst_n1678), .Y(aes_core_sbox_inst_n286) );
  NOR2X1 aes_core_sbox_inst_U748 ( .A(aes_core_sbox_inst_n46), .B(
        aes_core_sbox_inst_n35), .Y(aes_core_sbox_inst_n333) );
  AOI21X1 aes_core_sbox_inst_U747 ( .A0(aes_core_sbox_inst_n42), .A1(
        aes_core_sbox_inst_n87), .B0(aes_core_sbox_inst_n356), .Y(
        aes_core_sbox_inst_n311) );
  NOR2X1 aes_core_sbox_inst_U746 ( .A(aes_core_sbox_inst_n46), .B(
        aes_core_sbox_inst_n33), .Y(aes_core_sbox_inst_n1342) );
  OAI22X1 aes_core_sbox_inst_U745 ( .A0(aes_core_sbox_inst_n48), .A1(
        aes_core_sbox_inst_n1721), .B0(aes_core_sbox_inst_n186), .B1(
        aes_core_sbox_inst_n429), .Y(aes_core_sbox_inst_n428) );
  OAI22X1 aes_core_sbox_inst_U744 ( .A0(aes_core_sbox_inst_n21), .A1(
        aes_core_sbox_inst_n1603), .B0(aes_core_sbox_inst_n164), .B1(
        aes_core_sbox_inst_n1024), .Y(aes_core_sbox_inst_n1023) );
  OAI22X1 aes_core_sbox_inst_U743 ( .A0(aes_core_sbox_inst_n13), .A1(
        aes_core_sbox_inst_n244), .B0(aes_core_sbox_inst_n146), .B1(
        aes_core_sbox_inst_n662), .Y(aes_core_sbox_inst_n661) );
  OAI22X1 aes_core_sbox_inst_U742 ( .A0(aes_core_sbox_inst_n31), .A1(
        aes_core_sbox_inst_n1659), .B0(aes_core_sbox_inst_n179), .B1(
        aes_core_sbox_inst_n1362), .Y(aes_core_sbox_inst_n1361) );
  AOI21X1 aes_core_sbox_inst_U741 ( .A0(aes_core_sbox_inst_n194), .A1(
        aes_core_sbox_inst_n65), .B0(aes_core_sbox_inst_n68), .Y(
        aes_core_sbox_inst_n476) );
  AOI21X1 aes_core_sbox_inst_U740 ( .A0(aes_core_sbox_inst_n171), .A1(
        aes_core_sbox_inst_n91), .B0(aes_core_sbox_inst_n94), .Y(
        aes_core_sbox_inst_n1071) );
  AOI21X1 aes_core_sbox_inst_U739 ( .A0(aes_core_sbox_inst_n152), .A1(
        aes_core_sbox_inst_n105), .B0(aes_core_sbox_inst_n108), .Y(
        aes_core_sbox_inst_n709) );
  NOR2X1 aes_core_sbox_inst_U738 ( .A(aes_core_sbox_inst_n13), .B(
        aes_core_sbox_inst_n235), .Y(aes_core_sbox_inst_n947) );
  NOR2X1 aes_core_sbox_inst_U737 ( .A(aes_core_sbox_inst_n1725), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n430) );
  NOR2X1 aes_core_sbox_inst_U736 ( .A(aes_core_sbox_inst_n1607), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n1025) );
  NOR2X1 aes_core_sbox_inst_U735 ( .A(aes_core_sbox_inst_n248), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n663) );
  OAI211X1 aes_core_sbox_inst_U734 ( .A0(aes_core_sbox_inst_n19), .A1(
        aes_core_sbox_inst_n243), .B0(aes_core_sbox_inst_n662), .C0(
        aes_core_sbox_inst_n627), .Y(aes_core_sbox_inst_n762) );
  OAI211X1 aes_core_sbox_inst_U733 ( .A0(aes_core_sbox_inst_n81), .A1(
        aes_core_sbox_inst_n37), .B0(aes_core_sbox_inst_n1362), .C0(
        aes_core_sbox_inst_n1339), .Y(aes_core_sbox_inst_n1410) );
  AOI31X1 aes_core_sbox_inst_U732 ( .A0(aes_core_sbox_inst_n249), .A1(
        aes_core_sbox_inst_n248), .A2(aes_core_sbox_inst_n662), .B0(
        aes_core_sbox_inst_n215), .Y(aes_core_sbox_inst_n773) );
  INVX1 aes_core_sbox_inst_U731 ( .A(aes_core_sbox_inst_n592), .Y(
        aes_core_sbox_inst_n1684) );
  INVX1 aes_core_sbox_inst_U730 ( .A(aes_core_sbox_inst_n1217), .Y(
        aes_core_sbox_inst_n1566) );
  NOR2X1 aes_core_sbox_inst_U729 ( .A(aes_core_sbox_inst_n48), .B(
        aes_core_sbox_inst_n1703), .Y(aes_core_sbox_inst_n603) );
  NOR2X1 aes_core_sbox_inst_U728 ( .A(aes_core_sbox_inst_n21), .B(
        aes_core_sbox_inst_n22), .Y(aes_core_sbox_inst_n1228) );
  NOR2X1 aes_core_sbox_inst_U727 ( .A(aes_core_sbox_inst_n13), .B(
        aes_core_sbox_inst_n14), .Y(aes_core_sbox_inst_n870) );
  OAI22X1 aes_core_sbox_inst_U726 ( .A0(aes_core_sbox_inst_n221), .A1(
        aes_core_sbox_inst_n670), .B0(aes_core_sbox_inst_n118), .B1(
        aes_core_sbox_inst_n13), .Y(aes_core_sbox_inst_n668) );
  AOI221X1 aes_core_sbox_inst_U725 ( .A0(aes_core_sbox_inst_n15), .A1(
        aes_core_sbox_inst_n668), .B0(aes_core_sbox_inst_n108), .B1(
        aes_core_sbox_inst_n634), .C0(aes_core_sbox_inst_n669), .Y(
        aes_core_sbox_inst_n659) );
  NOR2X1 aes_core_sbox_inst_U724 ( .A(aes_core_sbox_inst_n36), .B(
        aes_core_sbox_inst_n81), .Y(aes_core_sbox_inst_n358) );
  AOI31X1 aes_core_sbox_inst_U723 ( .A0(aes_core_sbox_inst_n182), .A1(
        aes_core_sbox_inst_n47), .A2(aes_core_sbox_inst_n88), .B0(
        aes_core_sbox_inst_n288), .Y(aes_core_sbox_inst_n287) );
  NOR2X1 aes_core_sbox_inst_U722 ( .A(aes_core_sbox_inst_n237), .B(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n680) );
  AOI211X1 aes_core_sbox_inst_U721 ( .A0(aes_core_sbox_inst_n449), .A1(
        aes_core_sbox_inst_n192), .B0(aes_core_sbox_inst_n77), .C0(
        aes_core_sbox_inst_n422), .Y(aes_core_sbox_inst_n550) );
  AOI211X1 aes_core_sbox_inst_U720 ( .A0(aes_core_sbox_inst_n1044), .A1(
        aes_core_sbox_inst_n170), .B0(aes_core_sbox_inst_n103), .C0(
        aes_core_sbox_inst_n1017), .Y(aes_core_sbox_inst_n1145) );
  AOI211X1 aes_core_sbox_inst_U719 ( .A0(aes_core_sbox_inst_n682), .A1(
        aes_core_sbox_inst_n151), .B0(aes_core_sbox_inst_n115), .C0(
        aes_core_sbox_inst_n655), .Y(aes_core_sbox_inst_n817) );
  NOR3X1 aes_core_sbox_inst_U718 ( .A(aes_core_sbox_inst_n1691), .B(
        aes_core_sbox_inst_n138), .C(aes_core_sbox_inst_n1720), .Y(
        aes_core_sbox_inst_n400) );
  NOR3X1 aes_core_sbox_inst_U717 ( .A(aes_core_sbox_inst_n1573), .B(
        aes_core_sbox_inst_n129), .C(aes_core_sbox_inst_n24), .Y(
        aes_core_sbox_inst_n995) );
  NOR3X1 aes_core_sbox_inst_U716 ( .A(aes_core_sbox_inst_n215), .B(
        aes_core_sbox_inst_n134), .C(aes_core_sbox_inst_n243), .Y(
        aes_core_sbox_inst_n633) );
  NOR2X1 aes_core_sbox_inst_U715 ( .A(aes_core_sbox_inst_n248), .B(
        aes_core_sbox_inst_n215), .Y(aes_core_sbox_inst_n625) );
  NOR2X1 aes_core_sbox_inst_U714 ( .A(aes_core_sbox_inst_n1623), .B(
        aes_core_sbox_inst_n179), .Y(aes_core_sbox_inst_n265) );
  NOR2X1 aes_core_sbox_inst_U713 ( .A(aes_core_sbox_inst_n22), .B(
        aes_core_sbox_inst_n1573), .Y(aes_core_sbox_inst_n1019) );
  NOR2X1 aes_core_sbox_inst_U712 ( .A(aes_core_sbox_inst_n14), .B(
        aes_core_sbox_inst_n215), .Y(aes_core_sbox_inst_n657) );
  NOR2X1 aes_core_sbox_inst_U711 ( .A(aes_core_sbox_inst_n235), .B(
        aes_core_sbox_inst_n215), .Y(aes_core_sbox_inst_n686) );
  NOR2X1 aes_core_sbox_inst_U710 ( .A(aes_core_sbox_inst_n243), .B(
        aes_core_sbox_inst_n13), .Y(aes_core_sbox_inst_n656) );
  AOI222X1 aes_core_sbox_inst_U709 ( .A0(aes_core_sbox_inst_n87), .A1(
        aes_core_sbox_inst_n43), .B0(aes_core_sbox_inst_n88), .B1(
        aes_core_sbox_inst_n125), .C0(aes_core_sbox_inst_n81), .C1(
        aes_core_sbox_inst_n86), .Y(aes_core_sbox_inst_n1377) );
  NOR2X1 aes_core_sbox_inst_U708 ( .A(aes_core_sbox_inst_n255), .B(
        aes_core_sbox_inst_n147), .Y(aes_core_sbox_inst_n632) );
  NOR2X1 aes_core_sbox_inst_U707 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n49), .Y(aes_core_sbox_inst_n469) );
  NOR2X1 aes_core_sbox_inst_U706 ( .A(aes_core_sbox_inst_n27), .B(
        aes_core_sbox_inst_n23), .Y(aes_core_sbox_inst_n1064) );
  NOR2X1 aes_core_sbox_inst_U705 ( .A(aes_core_sbox_inst_n1720), .B(
        aes_core_sbox_inst_n51), .Y(aes_core_sbox_inst_n397) );
  BUFX3 aes_core_sbox_inst_U704 ( .A(aes_core_sbox_inst_n397), .Y(
        aes_core_sbox_inst_n72) );
  NOR2X1 aes_core_sbox_inst_U703 ( .A(aes_core_sbox_inst_n24), .B(
        aes_core_sbox_inst_n27), .Y(aes_core_sbox_inst_n992) );
  BUFX3 aes_core_sbox_inst_U702 ( .A(aes_core_sbox_inst_n992), .Y(
        aes_core_sbox_inst_n98) );
  NOR2X1 aes_core_sbox_inst_U701 ( .A(aes_core_sbox_inst_n39), .B(
        aes_core_sbox_inst_n37), .Y(aes_core_sbox_inst_n317) );
  BUFX3 aes_core_sbox_inst_U700 ( .A(aes_core_sbox_inst_n317), .Y(
        aes_core_sbox_inst_n86) );
  INVX1 aes_core_sbox_inst_U699 ( .A(aes_core_sbox_inst_n1103), .Y(
        aes_core_sbox_inst_n1608) );
  NAND4X1 aes_core_sbox_inst_U698 ( .A(aes_core_sbox_inst_n1412), .B(
        aes_core_sbox_inst_n1658), .C(aes_core_sbox_inst_n1649), .D(
        aes_core_sbox_inst_n320), .Y(aes_core_sbox_inst_n1430) );
  NAND4X1 aes_core_sbox_inst_U697 ( .A(aes_core_sbox_inst_n499), .B(
        aes_core_sbox_inst_n518), .C(aes_core_sbox_inst_n416), .D(
        aes_core_sbox_inst_n502), .Y(aes_core_sbox_inst_n516) );
  NAND4X1 aes_core_sbox_inst_U696 ( .A(aes_core_sbox_inst_n1094), .B(
        aes_core_sbox_inst_n1113), .C(aes_core_sbox_inst_n1011), .D(
        aes_core_sbox_inst_n1097), .Y(aes_core_sbox_inst_n1111) );
  NAND4X1 aes_core_sbox_inst_U695 ( .A(aes_core_sbox_inst_n766), .B(
        aes_core_sbox_inst_n785), .C(aes_core_sbox_inst_n649), .D(
        aes_core_sbox_inst_n769), .Y(aes_core_sbox_inst_n783) );
  NAND4X1 aes_core_sbox_inst_U694 ( .A(aes_core_sbox_inst_n395), .B(
        aes_core_sbox_inst_n1718), .C(aes_core_sbox_inst_n732), .D(
        aes_core_sbox_inst_n733), .Y(aes_core_sbox_inst_n731) );
  AOI22X1 aes_core_sbox_inst_U693 ( .A0(aes_core_sbox_inst_n186), .A1(
        aes_core_sbox_inst_n730), .B0(aes_core_sbox_inst_n731), .B1(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n728) );
  AOI221X1 aes_core_sbox_inst_U692 ( .A0(aes_core_sbox_inst_n392), .A1(
        aes_core_sbox_inst_n70), .B0(aes_core_sbox_inst_n424), .B1(
        aes_core_sbox_inst_n53), .C0(aes_core_sbox_inst_n425), .Y(
        aes_core_sbox_inst_n729) );
  AOI21X1 aes_core_sbox_inst_U691 ( .A0(aes_core_sbox_inst_n728), .A1(
        aes_core_sbox_inst_n729), .B0(aes_core_sbox_inst_n1680), .Y(
        aes_core_sbox_inst_n727) );
  NAND4X1 aes_core_sbox_inst_U690 ( .A(aes_core_sbox_inst_n990), .B(
        aes_core_sbox_inst_n1600), .C(aes_core_sbox_inst_n1237), .D(
        aes_core_sbox_inst_n1238), .Y(aes_core_sbox_inst_n1236) );
  AOI22X1 aes_core_sbox_inst_U689 ( .A0(aes_core_sbox_inst_n164), .A1(
        aes_core_sbox_inst_n1235), .B0(aes_core_sbox_inst_n1236), .B1(
        aes_core_sbox_inst_n166), .Y(aes_core_sbox_inst_n1233) );
  AOI221X1 aes_core_sbox_inst_U688 ( .A0(aes_core_sbox_inst_n987), .A1(
        aes_core_sbox_inst_n96), .B0(aes_core_sbox_inst_n1019), .B1(
        aes_core_sbox_inst_n29), .C0(aes_core_sbox_inst_n1020), .Y(
        aes_core_sbox_inst_n1234) );
  AOI21X1 aes_core_sbox_inst_U687 ( .A0(aes_core_sbox_inst_n1233), .A1(
        aes_core_sbox_inst_n1234), .B0(aes_core_sbox_inst_n273), .Y(
        aes_core_sbox_inst_n1232) );
  NAND4X1 aes_core_sbox_inst_U686 ( .A(aes_core_sbox_inst_n628), .B(
        aes_core_sbox_inst_n241), .C(aes_core_sbox_inst_n879), .D(
        aes_core_sbox_inst_n880), .Y(aes_core_sbox_inst_n878) );
  AOI22X1 aes_core_sbox_inst_U685 ( .A0(aes_core_sbox_inst_n146), .A1(
        aes_core_sbox_inst_n877), .B0(aes_core_sbox_inst_n878), .B1(
        aes_core_sbox_inst_n149), .Y(aes_core_sbox_inst_n875) );
  AOI221X1 aes_core_sbox_inst_U684 ( .A0(aes_core_sbox_inst_n625), .A1(
        aes_core_sbox_inst_n109), .B0(aes_core_sbox_inst_n657), .B1(
        aes_core_sbox_inst_n19), .C0(aes_core_sbox_inst_n658), .Y(
        aes_core_sbox_inst_n876) );
  AOI21X1 aes_core_sbox_inst_U683 ( .A0(aes_core_sbox_inst_n875), .A1(
        aes_core_sbox_inst_n876), .B0(aes_core_sbox_inst_n204), .Y(
        aes_core_sbox_inst_n874) );
  NAND4X1 aes_core_sbox_inst_U682 ( .A(aes_core_sbox_inst_n1639), .B(
        aes_core_sbox_inst_n1339), .C(aes_core_sbox_inst_n1666), .D(
        aes_core_sbox_inst_n319), .Y(aes_core_sbox_inst_n1453) );
  NOR2X1 aes_core_sbox_inst_U681 ( .A(aes_core_sbox_inst_n35), .B(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n282) );
  BUFX3 aes_core_sbox_inst_U680 ( .A(aes_core_sbox_inst_n282), .Y(
        aes_core_sbox_inst_n83) );
  NOR2X1 aes_core_sbox_inst_U679 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_sbox_inst_n22), .Y(aes_core_sbox_inst_n1057) );
  BUFX3 aes_core_sbox_inst_U678 ( .A(aes_core_sbox_inst_n1057), .Y(
        aes_core_sbox_inst_n101) );
  NOR2X1 aes_core_sbox_inst_U677 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n1703), .Y(aes_core_sbox_inst_n462) );
  BUFX3 aes_core_sbox_inst_U676 ( .A(aes_core_sbox_inst_n462), .Y(
        aes_core_sbox_inst_n75) );
  NOR2X1 aes_core_sbox_inst_U675 ( .A(aes_core_sbox_inst_n255), .B(
        aes_core_sbox_inst_n14), .Y(aes_core_sbox_inst_n695) );
  BUFX3 aes_core_sbox_inst_U674 ( .A(aes_core_sbox_inst_n695), .Y(
        aes_core_sbox_inst_n113) );
  CLKINVX3 aes_core_sbox_inst_U673 ( .A(aes_core_sbox_inst_n185), .Y(
        aes_core_sbox_inst_n179) );
  INVX1 aes_core_sbox_inst_U672 ( .A(aes_core_sbox_inst_n313), .Y(
        aes_core_sbox_inst_n1671) );
  AOI211X1 aes_core_sbox_inst_U671 ( .A0(aes_core_sbox_inst_n77), .A1(
        aes_core_sbox_inst_n53), .B0(aes_core_sbox_inst_n544), .C0(
        aes_core_sbox_inst_n524), .Y(aes_core_sbox_inst_n1181) );
  AOI22X1 aes_core_sbox_inst_U670 ( .A0(aes_core_sbox_inst_n75), .A1(
        aes_core_sbox_inst_n140), .B0(aes_core_sbox_inst_n138), .B1(
        aes_core_sbox_inst_n65), .Y(aes_core_sbox_inst_n1180) );
  AOI21X1 aes_core_sbox_inst_U669 ( .A0(aes_core_sbox_inst_n1180), .A1(
        aes_core_sbox_inst_n1181), .B0(aes_core_sbox_inst_n1683), .Y(
        aes_core_sbox_inst_n1175) );
  AOI211X1 aes_core_sbox_inst_U668 ( .A0(aes_core_sbox_inst_n103), .A1(
        aes_core_sbox_inst_n29), .B0(aes_core_sbox_inst_n1139), .C0(
        aes_core_sbox_inst_n1119), .Y(aes_core_sbox_inst_n1285) );
  AOI22X1 aes_core_sbox_inst_U667 ( .A0(aes_core_sbox_inst_n101), .A1(
        aes_core_sbox_inst_n133), .B0(aes_core_sbox_inst_n129), .B1(
        aes_core_sbox_inst_n91), .Y(aes_core_sbox_inst_n1284) );
  AOI21X1 aes_core_sbox_inst_U666 ( .A0(aes_core_sbox_inst_n1284), .A1(
        aes_core_sbox_inst_n1285), .B0(aes_core_sbox_inst_n617), .Y(
        aes_core_sbox_inst_n1279) );
  AOI211X1 aes_core_sbox_inst_U665 ( .A0(aes_core_sbox_inst_n115), .A1(
        aes_core_sbox_inst_n19), .B0(aes_core_sbox_inst_n811), .C0(
        aes_core_sbox_inst_n791), .Y(aes_core_sbox_inst_n927) );
  AOI22X1 aes_core_sbox_inst_U664 ( .A0(aes_core_sbox_inst_n113), .A1(
        aes_core_sbox_inst_n136), .B0(aes_core_sbox_inst_n134), .B1(
        aes_core_sbox_inst_n105), .Y(aes_core_sbox_inst_n926) );
  AOI21X1 aes_core_sbox_inst_U663 ( .A0(aes_core_sbox_inst_n926), .A1(
        aes_core_sbox_inst_n927), .B0(aes_core_sbox_inst_n207), .Y(
        aes_core_sbox_inst_n921) );
  NOR2X1 aes_core_sbox_inst_U662 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n1725), .Y(aes_core_sbox_inst_n484) );
  BUFX3 aes_core_sbox_inst_U661 ( .A(aes_core_sbox_inst_n484), .Y(
        aes_core_sbox_inst_n77) );
  NOR2X1 aes_core_sbox_inst_U660 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_sbox_inst_n1607), .Y(aes_core_sbox_inst_n1079) );
  BUFX3 aes_core_sbox_inst_U659 ( .A(aes_core_sbox_inst_n1079), .Y(
        aes_core_sbox_inst_n103) );
  NOR2X1 aes_core_sbox_inst_U658 ( .A(aes_core_sbox_inst_n18), .B(
        aes_core_sbox_inst_n248), .Y(aes_core_sbox_inst_n717) );
  BUFX3 aes_core_sbox_inst_U657 ( .A(aes_core_sbox_inst_n717), .Y(
        aes_core_sbox_inst_n115) );
  NAND2X1 aes_core_sbox_inst_U656 ( .A(aes_core_sbox_inst_n1724), .B(
        aes_core_sbox_inst_n1700), .Y(aes_core_sbox_inst_n381) );
  NAND2X1 aes_core_sbox_inst_U655 ( .A(aes_core_sbox_inst_n1606), .B(
        aes_core_sbox_inst_n1582), .Y(aes_core_sbox_inst_n976) );
  NAND2X1 aes_core_sbox_inst_U654 ( .A(aes_core_sbox_inst_n247), .B(
        aes_core_sbox_inst_n11), .Y(aes_core_sbox_inst_n614) );
  INVX1 aes_core_sbox_inst_U653 ( .A(aes_core_sbox_inst_n1356), .Y(
        aes_core_sbox_inst_n1650) );
  NAND2X1 aes_core_sbox_inst_U652 ( .A(aes_core_sbox_inst_n1661), .B(
        aes_core_sbox_inst_n1654), .Y(aes_core_sbox_inst_n1333) );
  OAI22X1 aes_core_sbox_inst_U651 ( .A0(aes_core_sbox_inst_n35), .A1(
        aes_core_sbox_inst_n42), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n32), .Y(aes_core_sbox_inst_n1437) );
  NAND2X1 aes_core_sbox_inst_U650 ( .A(aes_core_sbox_inst_n32), .B(
        aes_core_sbox_inst_n1664), .Y(aes_core_sbox_inst_n283) );
  NOR2X1 aes_core_sbox_inst_U649 ( .A(aes_core_sbox_inst_n48), .B(
        aes_core_sbox_inst_n1712), .Y(aes_core_sbox_inst_n1547) );
  NOR2X1 aes_core_sbox_inst_U648 ( .A(aes_core_sbox_inst_n21), .B(
        aes_core_sbox_inst_n1594), .Y(aes_core_sbox_inst_n1305) );
  AOI22X1 aes_core_sbox_inst_U647 ( .A0(aes_core_sbox_inst_n42), .A1(
        aes_core_sbox_inst_n88), .B0(aes_core_sbox_inst_n83), .B1(
        aes_core_sbox_inst_n81), .Y(aes_core_sbox_inst_n1364) );
  NAND2X1 aes_core_sbox_inst_U646 ( .A(aes_core_sbox_inst_n1709), .B(
        aes_core_sbox_inst_n1714), .Y(aes_core_sbox_inst_n742) );
  NAND2X1 aes_core_sbox_inst_U645 ( .A(aes_core_sbox_inst_n1591), .B(
        aes_core_sbox_inst_n1596), .Y(aes_core_sbox_inst_n1247) );
  NAND2X1 aes_core_sbox_inst_U644 ( .A(aes_core_sbox_inst_n232), .B(
        aes_core_sbox_inst_n237), .Y(aes_core_sbox_inst_n889) );
  OAI211X1 aes_core_sbox_inst_U643 ( .A0(aes_core_sbox_inst_n53), .A1(
        aes_core_sbox_inst_n1720), .B0(aes_core_sbox_inst_n429), .C0(
        aes_core_sbox_inst_n394), .Y(aes_core_sbox_inst_n495) );
  OAI211X1 aes_core_sbox_inst_U642 ( .A0(aes_core_sbox_inst_n29), .A1(
        aes_core_sbox_inst_n24), .B0(aes_core_sbox_inst_n1024), .C0(
        aes_core_sbox_inst_n989), .Y(aes_core_sbox_inst_n1090) );
  AOI31X1 aes_core_sbox_inst_U641 ( .A0(aes_core_sbox_inst_n1726), .A1(
        aes_core_sbox_inst_n1725), .A2(aes_core_sbox_inst_n429), .B0(
        aes_core_sbox_inst_n1691), .Y(aes_core_sbox_inst_n506) );
  AOI31X1 aes_core_sbox_inst_U640 ( .A0(aes_core_sbox_inst_n1608), .A1(
        aes_core_sbox_inst_n1607), .A2(aes_core_sbox_inst_n1024), .B0(
        aes_core_sbox_inst_n1573), .Y(aes_core_sbox_inst_n1101) );
  AOI31X1 aes_core_sbox_inst_U639 ( .A0(aes_core_sbox_inst_n1671), .A1(
        aes_core_sbox_inst_n35), .A2(aes_core_sbox_inst_n1362), .B0(
        aes_core_sbox_inst_n1630), .Y(aes_core_sbox_inst_n1420) );
  OAI211X1 aes_core_sbox_inst_U638 ( .A0(aes_core_sbox_inst_n44), .A1(
        aes_core_sbox_inst_n36), .B0(aes_core_sbox_inst_n319), .C0(
        aes_core_sbox_inst_n320), .Y(aes_core_sbox_inst_n318) );
  NAND2X1 aes_core_sbox_inst_U637 ( .A(aes_core_sbox_inst_n87), .B(
        aes_core_sbox_inst_n124), .Y(aes_core_sbox_inst_n337) );
  NOR2X1 aes_core_sbox_inst_U636 ( .A(aes_core_sbox_inst_n42), .B(
        aes_core_sbox_inst_n1660), .Y(aes_core_sbox_inst_n277) );
  AOI31X1 aes_core_sbox_inst_U635 ( .A0(aes_core_sbox_inst_n1721), .A1(
        aes_core_sbox_inst_n1705), .A2(aes_core_sbox_inst_n1699), .B0(
        aes_core_sbox_inst_n48), .Y(aes_core_sbox_inst_n414) );
  AOI31X1 aes_core_sbox_inst_U634 ( .A0(aes_core_sbox_inst_n1603), .A1(
        aes_core_sbox_inst_n1587), .A2(aes_core_sbox_inst_n1581), .B0(
        aes_core_sbox_inst_n21), .Y(aes_core_sbox_inst_n1009) );
  AOI31X1 aes_core_sbox_inst_U633 ( .A0(aes_core_sbox_inst_n244), .A1(
        aes_core_sbox_inst_n228), .A2(aes_core_sbox_inst_n223), .B0(
        aes_core_sbox_inst_n13), .Y(aes_core_sbox_inst_n647) );
  NOR2X1 aes_core_sbox_inst_U632 ( .A(aes_core_sbox_inst_n1723), .B(
        aes_core_sbox_inst_n194), .Y(aes_core_sbox_inst_n387) );
  NOR2X1 aes_core_sbox_inst_U631 ( .A(aes_core_sbox_inst_n1605), .B(
        aes_core_sbox_inst_n171), .Y(aes_core_sbox_inst_n982) );
  NOR2X1 aes_core_sbox_inst_U630 ( .A(aes_core_sbox_inst_n246), .B(
        aes_core_sbox_inst_n152), .Y(aes_core_sbox_inst_n620) );
  NOR2X1 aes_core_sbox_inst_U629 ( .A(aes_core_sbox_inst_n1664), .B(
        aes_core_sbox_inst_n124), .Y(aes_core_sbox_inst_n346) );
  AOI31X1 aes_core_sbox_inst_U628 ( .A0(aes_core_sbox_inst_n1659), .A1(
        aes_core_sbox_inst_n337), .A2(aes_core_sbox_inst_n1648), .B0(
        aes_core_sbox_inst_n31), .Y(aes_core_sbox_inst_n1352) );
  OAI22X1 aes_core_sbox_inst_U627 ( .A0(aes_core_sbox_inst_n1697), .A1(
        aes_core_sbox_inst_n69), .B0(aes_core_sbox_inst_n127), .B1(
        aes_core_sbox_inst_n48), .Y(aes_core_sbox_inst_n435) );
  AOI221X1 aes_core_sbox_inst_U626 ( .A0(aes_core_sbox_inst_n49), .A1(
        aes_core_sbox_inst_n435), .B0(aes_core_sbox_inst_n68), .B1(
        aes_core_sbox_inst_n401), .C0(aes_core_sbox_inst_n436), .Y(
        aes_core_sbox_inst_n426) );
  OAI22X1 aes_core_sbox_inst_U625 ( .A0(aes_core_sbox_inst_n1579), .A1(
        aes_core_sbox_inst_n95), .B0(aes_core_sbox_inst_n122), .B1(
        aes_core_sbox_inst_n21), .Y(aes_core_sbox_inst_n1030) );
  AOI221X1 aes_core_sbox_inst_U624 ( .A0(aes_core_sbox_inst_n23), .A1(
        aes_core_sbox_inst_n1030), .B0(aes_core_sbox_inst_n94), .B1(
        aes_core_sbox_inst_n996), .C0(aes_core_sbox_inst_n1031), .Y(
        aes_core_sbox_inst_n1021) );
  INVX1 aes_core_sbox_inst_U623 ( .A(aes_core_sbox_inst_n752), .Y(
        aes_core_sbox_inst_n1694) );
  AOI222X1 aes_core_sbox_inst_U622 ( .A0(aes_core_sbox_inst_n187), .A1(
        aes_core_sbox_inst_n1556), .B0(aes_core_sbox_inst_n1692), .B1(
        aes_core_sbox_inst_n128), .C0(aes_core_sbox_inst_n423), .C1(
        aes_core_sbox_inst_n54), .Y(aes_core_sbox_inst_n1555) );
  AOI31X1 aes_core_sbox_inst_U621 ( .A0(aes_core_sbox_inst_n70), .A1(
        aes_core_sbox_inst_n1704), .A2(aes_core_sbox_inst_n399), .B0(
        aes_core_sbox_inst_n1694), .Y(aes_core_sbox_inst_n1554) );
  OAI211X1 aes_core_sbox_inst_U620 ( .A0(aes_core_sbox_inst_n70), .A1(
        aes_core_sbox_inst_n1695), .B0(aes_core_sbox_inst_n1554), .C0(
        aes_core_sbox_inst_n1555), .Y(aes_core_sbox_inst_n1553) );
  INVX1 aes_core_sbox_inst_U619 ( .A(aes_core_sbox_inst_n1257), .Y(
        aes_core_sbox_inst_n1576) );
  AOI222X1 aes_core_sbox_inst_U618 ( .A0(aes_core_sbox_inst_n165), .A1(
        aes_core_sbox_inst_n1314), .B0(aes_core_sbox_inst_n1574), .B1(
        aes_core_sbox_inst_n123), .C0(aes_core_sbox_inst_n1018), .C1(
        aes_core_sbox_inst_n30), .Y(aes_core_sbox_inst_n1313) );
  AOI31X1 aes_core_sbox_inst_U617 ( .A0(aes_core_sbox_inst_n96), .A1(
        aes_core_sbox_inst_n1586), .A2(aes_core_sbox_inst_n994), .B0(
        aes_core_sbox_inst_n1576), .Y(aes_core_sbox_inst_n1312) );
  OAI211X1 aes_core_sbox_inst_U616 ( .A0(aes_core_sbox_inst_n96), .A1(
        aes_core_sbox_inst_n1577), .B0(aes_core_sbox_inst_n1312), .C0(
        aes_core_sbox_inst_n1313), .Y(aes_core_sbox_inst_n1311) );
  INVX1 aes_core_sbox_inst_U615 ( .A(aes_core_sbox_inst_n899), .Y(
        aes_core_sbox_inst_n218) );
  AOI222X1 aes_core_sbox_inst_U614 ( .A0(aes_core_sbox_inst_n147), .A1(
        aes_core_sbox_inst_n956), .B0(aes_core_sbox_inst_n216), .B1(
        aes_core_sbox_inst_n119), .C0(aes_core_sbox_inst_n656), .C1(
        aes_core_sbox_inst_n259), .Y(aes_core_sbox_inst_n955) );
  AOI31X1 aes_core_sbox_inst_U613 ( .A0(aes_core_sbox_inst_n109), .A1(
        aes_core_sbox_inst_n227), .A2(aes_core_sbox_inst_n632), .B0(
        aes_core_sbox_inst_n218), .Y(aes_core_sbox_inst_n954) );
  OAI211X1 aes_core_sbox_inst_U612 ( .A0(aes_core_sbox_inst_n109), .A1(
        aes_core_sbox_inst_n219), .B0(aes_core_sbox_inst_n954), .C0(
        aes_core_sbox_inst_n955), .Y(aes_core_sbox_inst_n953) );
  NOR2X1 aes_core_sbox_inst_U611 ( .A(aes_core_sbox_inst_n1714), .B(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n447) );
  NOR2X1 aes_core_sbox_inst_U610 ( .A(aes_core_sbox_inst_n1596), .B(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1042) );
  NAND4X1 aes_core_sbox_inst_U609 ( .A(aes_core_sbox_inst_n353), .B(
        aes_core_sbox_inst_n319), .C(aes_core_sbox_inst_n354), .D(
        aes_core_sbox_inst_n355), .Y(aes_core_sbox_inst_n351) );
  AOI31X1 aes_core_sbox_inst_U608 ( .A0(aes_core_sbox_inst_n1656), .A1(
        aes_core_sbox_inst_n125), .A2(aes_core_sbox_inst_n359), .B0(
        aes_core_sbox_inst_n1633), .Y(aes_core_sbox_inst_n349) );
  AOI222X1 aes_core_sbox_inst_U607 ( .A0(aes_core_sbox_inst_n179), .A1(
        aes_core_sbox_inst_n351), .B0(aes_core_sbox_inst_n1631), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n352), .C1(
        aes_core_sbox_inst_n1677), .Y(aes_core_sbox_inst_n350) );
  OAI211X1 aes_core_sbox_inst_U606 ( .A0(aes_core_sbox_inst_n125), .A1(
        aes_core_sbox_inst_n338), .B0(aes_core_sbox_inst_n349), .C0(
        aes_core_sbox_inst_n350), .Y(aes_core_sbox_inst_n348) );
  NOR2X1 aes_core_sbox_inst_U605 ( .A(aes_core_sbox_inst_n31), .B(
        aes_core_sbox_inst_n33), .Y(aes_core_sbox_inst_n1397) );
  NOR2X1 aes_core_sbox_inst_U604 ( .A(aes_core_sbox_inst_n1630), .B(
        aes_core_sbox_inst_n33), .Y(aes_core_sbox_inst_n290) );
  NAND2X1 aes_core_sbox_inst_U603 ( .A(aes_core_sbox_inst_n356), .B(
        aes_core_sbox_inst_n46), .Y(aes_core_sbox_inst_n1340) );
  NOR2X1 aes_core_sbox_inst_U602 ( .A(aes_core_sbox_inst_n31), .B(
        aes_core_sbox_inst_n37), .Y(aes_core_sbox_inst_n352) );
  NOR3X1 aes_core_sbox_inst_U601 ( .A(aes_core_sbox_inst_n37), .B(
        aes_core_sbox_inst_n143), .C(aes_core_sbox_inst_n1630), .Y(
        aes_core_sbox_inst_n1343) );
  OAI211X1 aes_core_sbox_inst_U600 ( .A0(aes_core_sbox_inst_n1661), .A1(
        aes_core_sbox_inst_n125), .B0(aes_core_sbox_inst_n1665), .C0(
        aes_core_sbox_inst_n1639), .Y(aes_core_sbox_inst_n306) );
  AOI221X1 aes_core_sbox_inst_U599 ( .A0(aes_core_sbox_inst_n88), .A1(
        aes_core_sbox_inst_n144), .B0(aes_core_sbox_inst_n143), .B1(
        aes_core_sbox_inst_n87), .C0(aes_core_sbox_inst_n306), .Y(
        aes_core_sbox_inst_n304) );
  INVX1 aes_core_sbox_inst_U598 ( .A(aes_core_sbox_inst_n307), .Y(
        aes_core_sbox_inst_n1629) );
  OAI32X1 aes_core_sbox_inst_U597 ( .A0(aes_core_sbox_inst_n1629), .A1(
        aes_core_sbox_inst_n143), .A2(aes_core_sbox_inst_n1623), .B0(
        aes_core_sbox_inst_n304), .B1(aes_core_sbox_inst_n1621), .Y(
        aes_core_sbox_inst_n298) );
  NOR2X1 aes_core_sbox_inst_U596 ( .A(aes_core_sbox_inst_n1712), .B(
        aes_core_sbox_inst_n1691), .Y(aes_core_sbox_inst_n453) );
  NOR2X1 aes_core_sbox_inst_U595 ( .A(aes_core_sbox_inst_n1594), .B(
        aes_core_sbox_inst_n1573), .Y(aes_core_sbox_inst_n1048) );
  NOR2X1 aes_core_sbox_inst_U594 ( .A(aes_core_sbox_inst_n1630), .B(
        aes_core_sbox_inst_n1645), .Y(aes_core_sbox_inst_n291) );
  NOR2X1 aes_core_sbox_inst_U593 ( .A(aes_core_sbox_inst_n1720), .B(
        aes_core_sbox_inst_n48), .Y(aes_core_sbox_inst_n423) );
  NOR2X1 aes_core_sbox_inst_U592 ( .A(aes_core_sbox_inst_n24), .B(
        aes_core_sbox_inst_n21), .Y(aes_core_sbox_inst_n1018) );
  INVX1 aes_core_sbox_inst_U591 ( .A(aes_core_sbox_inst_n87), .Y(
        aes_core_sbox_inst_n1645) );
  INVX1 aes_core_sbox_inst_U590 ( .A(aes_core_sbox_inst_n105), .Y(
        aes_core_sbox_inst_n235) );
  INVX1 aes_core_sbox_inst_U589 ( .A(aes_core_sbox_inst_n65), .Y(
        aes_core_sbox_inst_n1712) );
  INVX1 aes_core_sbox_inst_U588 ( .A(aes_core_sbox_inst_n195), .Y(
        aes_core_sbox_inst_n192) );
  INVX1 aes_core_sbox_inst_U587 ( .A(aes_core_sbox_inst_n172), .Y(
        aes_core_sbox_inst_n170) );
  INVX1 aes_core_sbox_inst_U586 ( .A(aes_core_sbox_inst_n631), .Y(
        aes_core_sbox_inst_n223) );
  INVX1 aes_core_sbox_inst_U585 ( .A(aes_core_sbox_inst_n263), .Y(
        aes_core_sbox_inst_n1621) );
  NAND2X1 aes_core_sbox_inst_U584 ( .A(aes_core_sbox_inst_n469), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n478) );
  NAND2X1 aes_core_sbox_inst_U583 ( .A(aes_core_sbox_inst_n1064), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1073) );
  NAND2X1 aes_core_sbox_inst_U582 ( .A(aes_core_sbox_inst_n702), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n711) );
  NAND2X1 aes_core_sbox_inst_U581 ( .A(aes_core_sbox_inst_n9), .B(
        aes_core_sbox_inst_n630), .Y(aes_core_sbox_inst_n650) );
  INVX1 aes_core_sbox_inst_U580 ( .A(aes_core_sbox_inst_n630), .Y(
        aes_core_sbox_inst_n241) );
  INVX1 aes_core_sbox_inst_U579 ( .A(aes_core_sbox_inst_n424), .Y(
        aes_core_sbox_inst_n1690) );
  INVX1 aes_core_sbox_inst_U578 ( .A(aes_core_sbox_inst_n1019), .Y(
        aes_core_sbox_inst_n1572) );
  INVX1 aes_core_sbox_inst_U577 ( .A(aes_core_sbox_inst_n190), .Y(
        aes_core_sbox_inst_n187) );
  INVX1 aes_core_sbox_inst_U576 ( .A(aes_core_sbox_inst_n168), .Y(
        aes_core_sbox_inst_n165) );
  INVX1 aes_core_sbox_inst_U575 ( .A(aes_core_sbox_inst_n149), .Y(
        aes_core_sbox_inst_n147) );
  CLKINVX3 aes_core_sbox_inst_U574 ( .A(aes_core_sbox_inst_n81), .Y(
        aes_core_sbox_inst_n125) );
  AOI21X1 aes_core_sbox_inst_U573 ( .A0(aes_core_sbox_inst_n657), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n658), .Y(
        aes_core_sbox_inst_n645) );
  INVX1 aes_core_sbox_inst_U572 ( .A(aes_core_sbox_inst_n398), .Y(
        aes_core_sbox_inst_n1699) );
  INVX1 aes_core_sbox_inst_U571 ( .A(aes_core_sbox_inst_n993), .Y(
        aes_core_sbox_inst_n1581) );
  AND2X2 aes_core_sbox_inst_U570 ( .A(aes_core_sbox_inst_n686), .B(
        aes_core_sbox_inst_n154), .Y(aes_core_sbox_inst_n658) );
  AOI21X1 aes_core_sbox_inst_U569 ( .A0(aes_core_sbox_inst_n32), .A1(
        aes_core_sbox_inst_n337), .B0(aes_core_sbox_inst_n179), .Y(
        aes_core_sbox_inst_n1480) );
  INVX1 aes_core_sbox_inst_U568 ( .A(aes_core_sbox_inst_n1342), .Y(
        aes_core_sbox_inst_n1648) );
  INVX1 aes_core_sbox_inst_U567 ( .A(aes_core_sbox_inst_n430), .Y(
        aes_core_sbox_inst_n1721) );
  INVX1 aes_core_sbox_inst_U566 ( .A(aes_core_sbox_inst_n1025), .Y(
        aes_core_sbox_inst_n1603) );
  INVX1 aes_core_sbox_inst_U565 ( .A(aes_core_sbox_inst_n663), .Y(
        aes_core_sbox_inst_n244) );
  AOI21X1 aes_core_sbox_inst_U564 ( .A0(aes_core_sbox_inst_n1704), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n69), .Y(
        aes_core_sbox_inst_n1543) );
  AOI21X1 aes_core_sbox_inst_U563 ( .A0(aes_core_sbox_inst_n1586), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n95), .Y(
        aes_core_sbox_inst_n1301) );
  AOI21X1 aes_core_sbox_inst_U562 ( .A0(aes_core_sbox_inst_n227), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n670), .Y(
        aes_core_sbox_inst_n943) );
  NAND2X1 aes_core_sbox_inst_U561 ( .A(aes_core_sbox_inst_n603), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n752) );
  NAND2X1 aes_core_sbox_inst_U560 ( .A(aes_core_sbox_inst_n1228), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n1257) );
  NAND2X1 aes_core_sbox_inst_U559 ( .A(aes_core_sbox_inst_n870), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n899) );
  NOR2X1 aes_core_sbox_inst_U558 ( .A(aes_core_sbox_inst_n1718), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n563) );
  NAND2X1 aes_core_sbox_inst_U557 ( .A(aes_core_sbox_inst_n115), .B(
        aes_core_sbox_inst_n8), .Y(aes_core_sbox_inst_n627) );
  NAND2X1 aes_core_sbox_inst_U556 ( .A(aes_core_sbox_inst_n5), .B(
        aes_core_sbox_inst_n72), .Y(aes_core_sbox_inst_n417) );
  NAND2X1 aes_core_sbox_inst_U555 ( .A(aes_core_sbox_inst_n4), .B(
        aes_core_sbox_inst_n98), .Y(aes_core_sbox_inst_n1012) );
  OAI22X1 aes_core_sbox_inst_U554 ( .A0(aes_core_sbox_inst_n1645), .A1(
        aes_core_sbox_inst_n44), .B0(aes_core_sbox_inst_n45), .B1(
        aes_core_sbox_inst_n1637), .Y(aes_core_sbox_inst_n1456) );
  OAI22X1 aes_core_sbox_inst_U553 ( .A0(aes_core_sbox_inst_n1712), .A1(
        aes_core_sbox_inst_n1735), .B0(aes_core_sbox_inst_n127), .B1(
        aes_core_sbox_inst_n1698), .Y(aes_core_sbox_inst_n546) );
  OAI22X1 aes_core_sbox_inst_U552 ( .A0(aes_core_sbox_inst_n1594), .A1(
        aes_core_sbox_inst_n1617), .B0(aes_core_sbox_inst_n122), .B1(
        aes_core_sbox_inst_n1580), .Y(aes_core_sbox_inst_n1141) );
  OAI22X1 aes_core_sbox_inst_U551 ( .A0(aes_core_sbox_inst_n235), .A1(
        aes_core_sbox_inst_n20), .B0(aes_core_sbox_inst_n118), .B1(
        aes_core_sbox_inst_n222), .Y(aes_core_sbox_inst_n813) );
  NAND2X1 aes_core_sbox_inst_U550 ( .A(aes_core_sbox_inst_n115), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n644) );
  AOI22X1 aes_core_sbox_inst_U549 ( .A0(aes_core_sbox_inst_n126), .A1(
        aes_core_sbox_inst_n77), .B0(aes_core_sbox_inst_n383), .B1(
        aes_core_sbox_inst_n469), .Y(aes_core_sbox_inst_n459) );
  AOI22X1 aes_core_sbox_inst_U548 ( .A0(aes_core_sbox_inst_n121), .A1(
        aes_core_sbox_inst_n103), .B0(aes_core_sbox_inst_n7), .B1(
        aes_core_sbox_inst_n1064), .Y(aes_core_sbox_inst_n1054) );
  AOI22X1 aes_core_sbox_inst_U547 ( .A0(aes_core_sbox_inst_n117), .A1(
        aes_core_sbox_inst_n115), .B0(aes_core_sbox_inst_n8), .B1(
        aes_core_sbox_inst_n702), .Y(aes_core_sbox_inst_n692) );
  INVX1 aes_core_sbox_inst_U546 ( .A(aes_core_sbox_inst_n399), .Y(
        aes_core_sbox_inst_n1697) );
  INVX1 aes_core_sbox_inst_U545 ( .A(aes_core_sbox_inst_n994), .Y(
        aes_core_sbox_inst_n1579) );
  NAND2X1 aes_core_sbox_inst_U544 ( .A(aes_core_sbox_inst_n75), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n416) );
  NAND2X1 aes_core_sbox_inst_U543 ( .A(aes_core_sbox_inst_n101), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n1011) );
  NAND2X1 aes_core_sbox_inst_U542 ( .A(aes_core_sbox_inst_n113), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n649) );
  INVX1 aes_core_sbox_inst_U541 ( .A(aes_core_sbox_inst_n359), .Y(
        aes_core_sbox_inst_n1636) );
  NOR2X1 aes_core_sbox_inst_U540 ( .A(aes_core_sbox_inst_n202), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n383) );
  NOR2X1 aes_core_sbox_inst_U539 ( .A(aes_core_sbox_inst_n177), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n978) );
  NOR2X1 aes_core_sbox_inst_U538 ( .A(aes_core_sbox_inst_n163), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n616) );
  NAND2X1 aes_core_sbox_inst_U537 ( .A(aes_core_sbox_inst_n67), .B(
        aes_core_sbox_inst_n75), .Y(aes_core_sbox_inst_n535) );
  NAND2X1 aes_core_sbox_inst_U536 ( .A(aes_core_sbox_inst_n93), .B(
        aes_core_sbox_inst_n101), .Y(aes_core_sbox_inst_n1130) );
  NAND2X1 aes_core_sbox_inst_U535 ( .A(aes_core_sbox_inst_n107), .B(
        aes_core_sbox_inst_n113), .Y(aes_core_sbox_inst_n802) );
  INVX1 aes_core_sbox_inst_U534 ( .A(aes_core_sbox_inst_n356), .Y(
        aes_core_sbox_inst_n1641) );
  BUFX3 aes_core_sbox_inst_U533 ( .A(aes_core_sbox_inst_n1641), .Y(
        aes_core_sbox_inst_n32) );
  INVX1 aes_core_sbox_inst_U532 ( .A(aes_core_sbox_inst_n395), .Y(
        aes_core_sbox_inst_n1711) );
  AOI21X1 aes_core_sbox_inst_U531 ( .A0(aes_core_sbox_inst_n127), .A1(
        aes_core_sbox_inst_n72), .B0(aes_core_sbox_inst_n1711), .Y(
        aes_core_sbox_inst_n432) );
  AOI21X1 aes_core_sbox_inst_U530 ( .A0(aes_core_sbox_inst_n424), .A1(
        aes_core_sbox_inst_n193), .B0(aes_core_sbox_inst_n425), .Y(
        aes_core_sbox_inst_n412) );
  AOI21X1 aes_core_sbox_inst_U529 ( .A0(aes_core_sbox_inst_n1019), .A1(
        aes_core_sbox_inst_n171), .B0(aes_core_sbox_inst_n1020), .Y(
        aes_core_sbox_inst_n1007) );
  AND2X2 aes_core_sbox_inst_U528 ( .A(aes_core_sbox_inst_n453), .B(
        aes_core_sbox_inst_n192), .Y(aes_core_sbox_inst_n425) );
  AND2X2 aes_core_sbox_inst_U527 ( .A(aes_core_sbox_inst_n1048), .B(
        aes_core_sbox_inst_n170), .Y(aes_core_sbox_inst_n1020) );
  CLKINVX3 aes_core_sbox_inst_U526 ( .A(aes_core_sbox_inst_n302), .Y(
        aes_core_sbox_inst_n124) );
  INVX1 aes_core_sbox_inst_U525 ( .A(aes_core_sbox_inst_n334), .Y(
        aes_core_sbox_inst_n1639) );
  CLKINVX3 aes_core_sbox_inst_U524 ( .A(aes_core_sbox_inst_n190), .Y(
        aes_core_sbox_inst_n186) );
  CLKINVX3 aes_core_sbox_inst_U523 ( .A(aes_core_sbox_inst_n168), .Y(
        aes_core_sbox_inst_n164) );
  NOR2X1 aes_core_sbox_inst_U522 ( .A(aes_core_sbox_inst_n194), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n472) );
  BUFX3 aes_core_sbox_inst_U521 ( .A(aes_core_sbox_inst_n472), .Y(
        aes_core_sbox_inst_n67) );
  NOR2X1 aes_core_sbox_inst_U520 ( .A(aes_core_sbox_inst_n173), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1067) );
  BUFX3 aes_core_sbox_inst_U519 ( .A(aes_core_sbox_inst_n1067), .Y(
        aes_core_sbox_inst_n93) );
  NAND2X1 aes_core_sbox_inst_U518 ( .A(aes_core_sbox_inst_n1397), .B(
        aes_core_sbox_inst_n40), .Y(aes_core_sbox_inst_n370) );
  INVX1 aes_core_sbox_inst_U517 ( .A(aes_core_sbox_inst_n1355), .Y(
        aes_core_sbox_inst_n1649) );
  CLKINVX3 aes_core_sbox_inst_U516 ( .A(aes_core_sbox_inst_n172), .Y(
        aes_core_sbox_inst_n169) );
  CLKINVX3 aes_core_sbox_inst_U515 ( .A(aes_core_sbox_inst_n195), .Y(
        aes_core_sbox_inst_n191) );
  CLKINVX3 aes_core_sbox_inst_U514 ( .A(aes_core_sbox_inst_n153), .Y(
        aes_core_sbox_inst_n151) );
  NOR2X1 aes_core_sbox_inst_U513 ( .A(aes_core_sbox_inst_n153), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n705) );
  BUFX3 aes_core_sbox_inst_U512 ( .A(aes_core_sbox_inst_n705), .Y(
        aes_core_sbox_inst_n107) );
  OAI22X1 aes_core_sbox_inst_U511 ( .A0(aes_core_sbox_inst_n138), .A1(
        aes_core_sbox_inst_n1709), .B0(aes_core_sbox_inst_n200), .B1(
        aes_core_sbox_inst_n1702), .Y(aes_core_sbox_inst_n1172) );
  AOI22X1 aes_core_sbox_inst_U510 ( .A0(aes_core_sbox_inst_n186), .A1(
        aes_core_sbox_inst_n1172), .B0(aes_core_sbox_inst_n424), .B1(
        aes_core_sbox_inst_n127), .Y(aes_core_sbox_inst_n1170) );
  OAI22X1 aes_core_sbox_inst_U509 ( .A0(aes_core_sbox_inst_n129), .A1(
        aes_core_sbox_inst_n1591), .B0(aes_core_sbox_inst_n177), .B1(
        aes_core_sbox_inst_n1584), .Y(aes_core_sbox_inst_n1276) );
  AOI22X1 aes_core_sbox_inst_U508 ( .A0(aes_core_sbox_inst_n164), .A1(
        aes_core_sbox_inst_n1276), .B0(aes_core_sbox_inst_n1019), .B1(
        aes_core_sbox_inst_n122), .Y(aes_core_sbox_inst_n1274) );
  OAI22X1 aes_core_sbox_inst_U507 ( .A0(aes_core_sbox_inst_n134), .A1(
        aes_core_sbox_inst_n232), .B0(aes_core_sbox_inst_n161), .B1(
        aes_core_sbox_inst_n225), .Y(aes_core_sbox_inst_n918) );
  AOI22X1 aes_core_sbox_inst_U506 ( .A0(aes_core_sbox_inst_n146), .A1(
        aes_core_sbox_inst_n918), .B0(aes_core_sbox_inst_n657), .B1(
        aes_core_sbox_inst_n118), .Y(aes_core_sbox_inst_n916) );
  NOR2X1 aes_core_sbox_inst_U505 ( .A(aes_core_sbox_inst_n40), .B(
        aes_core_sbox_inst_n36), .Y(aes_core_sbox_inst_n1432) );
  INVX1 aes_core_sbox_inst_U504 ( .A(aes_core_sbox_inst_n1528), .Y(
        aes_core_sbox_inst_n1640) );
  NAND2X1 aes_core_sbox_inst_U503 ( .A(aes_core_sbox_inst_n77), .B(
        aes_core_sbox_inst_n6), .Y(aes_core_sbox_inst_n394) );
  NAND2X1 aes_core_sbox_inst_U502 ( .A(aes_core_sbox_inst_n103), .B(
        aes_core_sbox_inst_n7), .Y(aes_core_sbox_inst_n989) );
  INVX1 aes_core_sbox_inst_U501 ( .A(aes_core_sbox_inst_n990), .Y(
        aes_core_sbox_inst_n1593) );
  AOI21X1 aes_core_sbox_inst_U500 ( .A0(aes_core_sbox_inst_n122), .A1(
        aes_core_sbox_inst_n98), .B0(aes_core_sbox_inst_n1593), .Y(
        aes_core_sbox_inst_n1027) );
  INVX1 aes_core_sbox_inst_U499 ( .A(aes_core_sbox_inst_n1340), .Y(
        aes_core_sbox_inst_n1642) );
  AOI21X1 aes_core_sbox_inst_U498 ( .A0(aes_core_sbox_inst_n1678), .A1(
        aes_core_sbox_inst_n86), .B0(aes_core_sbox_inst_n1642), .Y(
        aes_core_sbox_inst_n1365) );
  NOR2X1 aes_core_sbox_inst_U497 ( .A(aes_core_sbox_inst_n1661), .B(
        aes_core_sbox_inst_n179), .Y(aes_core_sbox_inst_n288) );
  NAND2X1 aes_core_sbox_inst_U496 ( .A(aes_core_sbox_inst_n77), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n411) );
  NAND2X1 aes_core_sbox_inst_U495 ( .A(aes_core_sbox_inst_n103), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n1006) );
  NOR2X1 aes_core_sbox_inst_U494 ( .A(aes_core_sbox_inst_n52), .B(
        aes_core_sbox_inst_n1712), .Y(aes_core_sbox_inst_n576) );
  NOR2X1 aes_core_sbox_inst_U493 ( .A(aes_core_sbox_inst_n28), .B(
        aes_core_sbox_inst_n1594), .Y(aes_core_sbox_inst_n1201) );
  AOI21X1 aes_core_sbox_inst_U492 ( .A0(aes_core_sbox_inst_n72), .A1(
        aes_core_sbox_inst_n191), .B0(aes_core_sbox_inst_n398), .Y(
        aes_core_sbox_inst_n396) );
  AOI31X1 aes_core_sbox_inst_U491 ( .A0(aes_core_sbox_inst_n394), .A1(
        aes_core_sbox_inst_n395), .A2(aes_core_sbox_inst_n396), .B0(
        aes_core_sbox_inst_n190), .Y(aes_core_sbox_inst_n393) );
  AOI21X1 aes_core_sbox_inst_U490 ( .A0(aes_core_sbox_inst_n98), .A1(
        aes_core_sbox_inst_n169), .B0(aes_core_sbox_inst_n993), .Y(
        aes_core_sbox_inst_n991) );
  AOI31X1 aes_core_sbox_inst_U489 ( .A0(aes_core_sbox_inst_n989), .A1(
        aes_core_sbox_inst_n990), .A2(aes_core_sbox_inst_n991), .B0(
        aes_core_sbox_inst_n168), .Y(aes_core_sbox_inst_n988) );
  AOI21X1 aes_core_sbox_inst_U488 ( .A0(aes_core_sbox_inst_n630), .A1(
        aes_core_sbox_inst_n151), .B0(aes_core_sbox_inst_n631), .Y(
        aes_core_sbox_inst_n629) );
  AOI31X1 aes_core_sbox_inst_U487 ( .A0(aes_core_sbox_inst_n627), .A1(
        aes_core_sbox_inst_n628), .A2(aes_core_sbox_inst_n629), .B0(
        aes_core_sbox_inst_n149), .Y(aes_core_sbox_inst_n626) );
  NOR2X1 aes_core_sbox_inst_U486 ( .A(aes_core_sbox_inst_n1709), .B(
        aes_core_sbox_inst_n200), .Y(aes_core_sbox_inst_n470) );
  NOR2X1 aes_core_sbox_inst_U485 ( .A(aes_core_sbox_inst_n1591), .B(
        aes_core_sbox_inst_n175), .Y(aes_core_sbox_inst_n1065) );
  NOR2X1 aes_core_sbox_inst_U484 ( .A(aes_core_sbox_inst_n232), .B(
        aes_core_sbox_inst_n163), .Y(aes_core_sbox_inst_n703) );
  INVX1 aes_core_sbox_inst_U483 ( .A(aes_core_sbox_inst_n1498), .Y(
        aes_core_sbox_inst_n1653) );
  AOI22X1 aes_core_sbox_inst_U482 ( .A0(aes_core_sbox_inst_n191), .A1(
        aes_core_sbox_inst_n72), .B0(aes_core_sbox_inst_n126), .B1(
        aes_core_sbox_inst_n77), .Y(aes_core_sbox_inst_n735) );
  AOI22X1 aes_core_sbox_inst_U481 ( .A0(aes_core_sbox_inst_n169), .A1(
        aes_core_sbox_inst_n98), .B0(aes_core_sbox_inst_n121), .B1(
        aes_core_sbox_inst_n103), .Y(aes_core_sbox_inst_n1240) );
  AOI22X1 aes_core_sbox_inst_U480 ( .A0(aes_core_sbox_inst_n151), .A1(
        aes_core_sbox_inst_n630), .B0(aes_core_sbox_inst_n117), .B1(
        aes_core_sbox_inst_n115), .Y(aes_core_sbox_inst_n882) );
  AOI22X1 aes_core_sbox_inst_U479 ( .A0(aes_core_sbox_inst_n193), .A1(
        aes_core_sbox_inst_n75), .B0(aes_core_sbox_inst_n52), .B1(
        aes_core_sbox_inst_n77), .Y(aes_core_sbox_inst_n431) );
  AOI22X1 aes_core_sbox_inst_U478 ( .A0(aes_core_sbox_inst_n171), .A1(
        aes_core_sbox_inst_n101), .B0(aes_core_sbox_inst_n28), .B1(
        aes_core_sbox_inst_n103), .Y(aes_core_sbox_inst_n1026) );
  AOI22X1 aes_core_sbox_inst_U477 ( .A0(aes_core_sbox_inst_n155), .A1(
        aes_core_sbox_inst_n113), .B0(aes_core_sbox_inst_n19), .B1(
        aes_core_sbox_inst_n115), .Y(aes_core_sbox_inst_n664) );
  AOI211X1 aes_core_sbox_inst_U476 ( .A0(aes_core_sbox_inst_n381), .A1(
        aes_core_sbox_inst_n54), .B0(aes_core_sbox_inst_n421), .C0(
        aes_core_sbox_inst_n602), .Y(aes_core_sbox_inst_n601) );
  AOI211X1 aes_core_sbox_inst_U475 ( .A0(aes_core_sbox_inst_n976), .A1(
        aes_core_sbox_inst_n30), .B0(aes_core_sbox_inst_n1016), .C0(
        aes_core_sbox_inst_n1227), .Y(aes_core_sbox_inst_n1226) );
  NOR2X1 aes_core_sbox_inst_U474 ( .A(aes_core_sbox_inst_n1709), .B(
        aes_core_sbox_inst_n194), .Y(aes_core_sbox_inst_n544) );
  NOR2X1 aes_core_sbox_inst_U473 ( .A(aes_core_sbox_inst_n1591), .B(
        aes_core_sbox_inst_n173), .Y(aes_core_sbox_inst_n1139) );
  NOR2X1 aes_core_sbox_inst_U472 ( .A(aes_core_sbox_inst_n232), .B(
        aes_core_sbox_inst_n152), .Y(aes_core_sbox_inst_n811) );
  NAND2X1 aes_core_sbox_inst_U471 ( .A(aes_core_sbox_inst_n68), .B(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n502) );
  NAND2X1 aes_core_sbox_inst_U470 ( .A(aes_core_sbox_inst_n94), .B(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1097) );
  NAND2X1 aes_core_sbox_inst_U469 ( .A(aes_core_sbox_inst_n108), .B(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n769) );
  AOI221X1 aes_core_sbox_inst_U468 ( .A0(aes_core_sbox_inst_n72), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n77), .B1(
        aes_core_sbox_inst_n128), .C0(aes_core_sbox_inst_n544), .Y(
        aes_core_sbox_inst_n1544) );
  AOI221X1 aes_core_sbox_inst_U467 ( .A0(aes_core_sbox_inst_n98), .A1(
        aes_core_sbox_inst_n121), .B0(aes_core_sbox_inst_n103), .B1(
        aes_core_sbox_inst_n123), .C0(aes_core_sbox_inst_n1139), .Y(
        aes_core_sbox_inst_n1302) );
  AOI221X1 aes_core_sbox_inst_U466 ( .A0(aes_core_sbox_inst_n630), .A1(
        aes_core_sbox_inst_n117), .B0(aes_core_sbox_inst_n115), .B1(
        aes_core_sbox_inst_n119), .C0(aes_core_sbox_inst_n811), .Y(
        aes_core_sbox_inst_n944) );
  AOI221X1 aes_core_sbox_inst_U465 ( .A0(aes_core_sbox_inst_n86), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n83), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n334), .Y(
        aes_core_sbox_inst_n331) );
  INVX1 aes_core_sbox_inst_U464 ( .A(aes_core_sbox_inst_n88), .Y(
        aes_core_sbox_inst_n1651) );
  INVX1 aes_core_sbox_inst_U463 ( .A(aes_core_sbox_inst_n108), .Y(
        aes_core_sbox_inst_n232) );
  INVX1 aes_core_sbox_inst_U462 ( .A(aes_core_sbox_inst_n68), .Y(
        aes_core_sbox_inst_n1709) );
  INVX1 aes_core_sbox_inst_U461 ( .A(aes_core_sbox_inst_n94), .Y(
        aes_core_sbox_inst_n1591) );
  NOR2X1 aes_core_sbox_inst_U460 ( .A(aes_core_sbox_inst_n107), .B(
        aes_core_sbox_inst_n146), .Y(aes_core_sbox_inst_n634) );
  INVX1 aes_core_sbox_inst_U459 ( .A(aes_core_sbox_inst_n670), .Y(
        aes_core_sbox_inst_n258) );
  INVX1 aes_core_sbox_inst_U458 ( .A(aes_core_sbox_inst_n258), .Y(
        aes_core_sbox_inst_n120) );
  INVX1 aes_core_sbox_inst_U457 ( .A(aes_core_sbox_inst_n384), .Y(
        aes_core_sbox_inst_n137) );
  INVX1 aes_core_sbox_inst_U456 ( .A(aes_core_sbox_inst_n142), .Y(
        aes_core_sbox_inst_n144) );
  INVX1 aes_core_sbox_inst_U455 ( .A(aes_core_sbox_inst_n383), .Y(
        aes_core_sbox_inst_n1735) );
  INVX1 aes_core_sbox_inst_U454 ( .A(aes_core_sbox_inst_n978), .Y(
        aes_core_sbox_inst_n1617) );
  INVX1 aes_core_sbox_inst_U453 ( .A(aes_core_sbox_inst_n616), .Y(
        aes_core_sbox_inst_n259) );
  INVX1 aes_core_sbox_inst_U452 ( .A(aes_core_sbox_inst_n1158), .Y(
        aes_core_sbox_inst_n1598) );
  INVX1 aes_core_sbox_inst_U451 ( .A(aes_core_sbox_inst_n830), .Y(
        aes_core_sbox_inst_n239) );
  NOR2X1 aes_core_sbox_inst_U450 ( .A(aes_core_sbox_inst_n219), .B(
        aes_core_sbox_inst_n136), .Y(aes_core_sbox_inst_n669) );
  OAI22X1 aes_core_sbox_inst_U449 ( .A0(aes_core_sbox_inst_n191), .A1(
        aes_core_sbox_inst_n1718), .B0(aes_core_sbox_inst_n1702), .B1(
        aes_core_sbox_inst_n127), .Y(aes_core_sbox_inst_n1551) );
  OAI22X1 aes_core_sbox_inst_U448 ( .A0(aes_core_sbox_inst_n151), .A1(
        aes_core_sbox_inst_n16), .B0(aes_core_sbox_inst_n225), .B1(
        aes_core_sbox_inst_n118), .Y(aes_core_sbox_inst_n951) );
  NOR2X1 aes_core_sbox_inst_U447 ( .A(aes_core_sbox_inst_n67), .B(
        aes_core_sbox_inst_n186), .Y(aes_core_sbox_inst_n401) );
  NOR2X1 aes_core_sbox_inst_U446 ( .A(aes_core_sbox_inst_n93), .B(
        aes_core_sbox_inst_n164), .Y(aes_core_sbox_inst_n996) );
  INVX1 aes_core_sbox_inst_U445 ( .A(aes_core_sbox_inst_n2), .Y(
        aes_core_sbox_inst_n142) );
  NAND2BX1 aes_core_sbox_inst_U444 ( .AN(aes_core_sbox_inst_n477), .B(
        aes_core_sbox_inst_n478), .Y(aes_core_sbox_inst_n475) );
  NAND2BX1 aes_core_sbox_inst_U443 ( .AN(aes_core_sbox_inst_n1072), .B(
        aes_core_sbox_inst_n1073), .Y(aes_core_sbox_inst_n1070) );
  NAND2BX1 aes_core_sbox_inst_U442 ( .AN(aes_core_sbox_inst_n710), .B(
        aes_core_sbox_inst_n711), .Y(aes_core_sbox_inst_n708) );
  NAND4BX1 aes_core_sbox_inst_U441 ( .AN(aes_core_sbox_inst_n544), .B(
        aes_core_sbox_inst_n394), .C(aes_core_sbox_inst_n1716), .D(
        aes_core_sbox_inst_n535), .Y(aes_core_sbox_inst_n542) );
  NAND4BX1 aes_core_sbox_inst_U440 ( .AN(aes_core_sbox_inst_n811), .B(
        aes_core_sbox_inst_n627), .C(aes_core_sbox_inst_n239), .D(
        aes_core_sbox_inst_n802), .Y(aes_core_sbox_inst_n809) );
  NOR2X1 aes_core_sbox_inst_U439 ( .A(aes_core_sbox_inst_n1695), .B(
        aes_core_sbox_inst_n140), .Y(aes_core_sbox_inst_n436) );
  NOR2X1 aes_core_sbox_inst_U438 ( .A(aes_core_sbox_inst_n1577), .B(
        aes_core_sbox_inst_n131), .Y(aes_core_sbox_inst_n1031) );
  NOR2X1 aes_core_sbox_inst_U437 ( .A(aes_core_sbox_inst_n1724), .B(
        aes_core_sbox_inst_n186), .Y(aes_core_sbox_inst_n405) );
  NOR2X1 aes_core_sbox_inst_U436 ( .A(aes_core_sbox_inst_n1606), .B(
        aes_core_sbox_inst_n164), .Y(aes_core_sbox_inst_n1000) );
  NOR2X1 aes_core_sbox_inst_U435 ( .A(aes_core_sbox_inst_n247), .B(
        aes_core_sbox_inst_n146), .Y(aes_core_sbox_inst_n638) );
  INVX1 aes_core_sbox_inst_U434 ( .A(aes_core_sbox_inst_n843), .Y(
        aes_core_sbox_inst_n228) );
  OAI22X1 aes_core_sbox_inst_U433 ( .A0(aes_core_sbox_inst_n169), .A1(
        aes_core_sbox_inst_n1600), .B0(aes_core_sbox_inst_n1584), .B1(
        aes_core_sbox_inst_n122), .Y(aes_core_sbox_inst_n1309) );
  NOR2X1 aes_core_sbox_inst_U432 ( .A(aes_core_sbox_inst_n232), .B(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n718) );
  AOI31X1 aes_core_sbox_inst_U431 ( .A0(aes_core_sbox_inst_n231), .A1(
        aes_core_sbox_inst_n649), .A2(aes_core_sbox_inst_n650), .B0(
        aes_core_sbox_inst_n147), .Y(aes_core_sbox_inst_n648) );
  NOR2X1 aes_core_sbox_inst_U430 ( .A(aes_core_sbox_inst_n1702), .B(
        aes_core_sbox_inst_n67), .Y(aes_core_sbox_inst_n422) );
  NOR2X1 aes_core_sbox_inst_U429 ( .A(aes_core_sbox_inst_n1584), .B(
        aes_core_sbox_inst_n93), .Y(aes_core_sbox_inst_n1017) );
  NOR2X1 aes_core_sbox_inst_U428 ( .A(aes_core_sbox_inst_n225), .B(
        aes_core_sbox_inst_n107), .Y(aes_core_sbox_inst_n655) );
  NOR2X1 aes_core_sbox_inst_U427 ( .A(aes_core_sbox_inst_n1702), .B(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n511) );
  NOR2X1 aes_core_sbox_inst_U426 ( .A(aes_core_sbox_inst_n1584), .B(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1106) );
  NOR2X1 aes_core_sbox_inst_U425 ( .A(aes_core_sbox_inst_n225), .B(
        aes_core_sbox_inst_n109), .Y(aes_core_sbox_inst_n778) );
  OAI211X1 aes_core_sbox_inst_U424 ( .A0(aes_core_sbox_inst_n192), .A1(
        aes_core_sbox_inst_n1702), .B0(aes_core_sbox_inst_n1707), .C0(
        aes_core_sbox_inst_n735), .Y(aes_core_sbox_inst_n730) );
  OAI211X1 aes_core_sbox_inst_U423 ( .A0(aes_core_sbox_inst_n170), .A1(
        aes_core_sbox_inst_n1584), .B0(aes_core_sbox_inst_n1589), .C0(
        aes_core_sbox_inst_n1240), .Y(aes_core_sbox_inst_n1235) );
  OAI211X1 aes_core_sbox_inst_U422 ( .A0(aes_core_sbox_inst_n154), .A1(
        aes_core_sbox_inst_n225), .B0(aes_core_sbox_inst_n230), .C0(
        aes_core_sbox_inst_n882), .Y(aes_core_sbox_inst_n877) );
  NOR2X1 aes_core_sbox_inst_U421 ( .A(aes_core_sbox_inst_n1709), .B(
        aes_core_sbox_inst_n70), .Y(aes_core_sbox_inst_n485) );
  NOR2X1 aes_core_sbox_inst_U420 ( .A(aes_core_sbox_inst_n1591), .B(
        aes_core_sbox_inst_n96), .Y(aes_core_sbox_inst_n1080) );
  AOI31X1 aes_core_sbox_inst_U419 ( .A0(aes_core_sbox_inst_n1708), .A1(
        aes_core_sbox_inst_n416), .A2(aes_core_sbox_inst_n417), .B0(
        aes_core_sbox_inst_n187), .Y(aes_core_sbox_inst_n415) );
  AOI31X1 aes_core_sbox_inst_U418 ( .A0(aes_core_sbox_inst_n1590), .A1(
        aes_core_sbox_inst_n1011), .A2(aes_core_sbox_inst_n1012), .B0(
        aes_core_sbox_inst_n165), .Y(aes_core_sbox_inst_n1010) );
  NOR2X1 aes_core_sbox_inst_U417 ( .A(aes_core_sbox_inst_n126), .B(
        aes_core_sbox_inst_n1709), .Y(aes_core_sbox_inst_n421) );
  NOR2X1 aes_core_sbox_inst_U416 ( .A(aes_core_sbox_inst_n121), .B(
        aes_core_sbox_inst_n1591), .Y(aes_core_sbox_inst_n1016) );
  INVX1 aes_core_sbox_inst_U415 ( .A(aes_core_sbox_inst_n135), .Y(
        aes_core_sbox_inst_n136) );
  INVX1 aes_core_sbox_inst_U414 ( .A(aes_core_sbox_inst_n1425), .Y(
        aes_core_sbox_inst_n1668) );
  INVX1 aes_core_sbox_inst_U413 ( .A(aes_core_sbox_inst_n655), .Y(
        aes_core_sbox_inst_n224) );
  NOR2X1 aes_core_sbox_inst_U412 ( .A(aes_core_sbox_inst_n16), .B(
        aes_core_sbox_inst_n134), .Y(aes_core_sbox_inst_n869) );
  INVX1 aes_core_sbox_inst_U411 ( .A(aes_core_sbox_inst_n142), .Y(
        aes_core_sbox_inst_n145) );
  INVX1 aes_core_sbox_inst_U410 ( .A(aes_core_sbox_inst_n70), .Y(
        aes_core_sbox_inst_n1734) );
  INVX1 aes_core_sbox_inst_U409 ( .A(aes_core_sbox_inst_n96), .Y(
        aes_core_sbox_inst_n1616) );
  INVX1 aes_core_sbox_inst_U408 ( .A(aes_core_sbox_inst_n109), .Y(
        aes_core_sbox_inst_n257) );
  CLKINVX3 aes_core_sbox_inst_U407 ( .A(aes_core_sbox_inst_n472), .Y(
        aes_core_sbox_inst_n126) );
  CLKINVX3 aes_core_sbox_inst_U406 ( .A(aes_core_sbox_inst_n1067), .Y(
        aes_core_sbox_inst_n121) );
  CLKINVX3 aes_core_sbox_inst_U405 ( .A(aes_core_sbox_inst_n705), .Y(
        aes_core_sbox_inst_n117) );
  INVX1 aes_core_sbox_inst_U404 ( .A(aes_core_sbox_inst_n422), .Y(
        aes_core_sbox_inst_n1701) );
  INVX1 aes_core_sbox_inst_U403 ( .A(aes_core_sbox_inst_n1017), .Y(
        aes_core_sbox_inst_n1583) );
  NOR2X1 aes_core_sbox_inst_U402 ( .A(aes_core_sbox_inst_n1718), .B(
        aes_core_sbox_inst_n138), .Y(aes_core_sbox_inst_n602) );
  NOR2X1 aes_core_sbox_inst_U401 ( .A(aes_core_sbox_inst_n1600), .B(
        aes_core_sbox_inst_n129), .Y(aes_core_sbox_inst_n1227) );
  INVX1 aes_core_sbox_inst_U400 ( .A(aes_core_sbox_inst_n485), .Y(
        aes_core_sbox_inst_n1708) );
  INVX1 aes_core_sbox_inst_U399 ( .A(aes_core_sbox_inst_n1080), .Y(
        aes_core_sbox_inst_n1590) );
  INVX1 aes_core_sbox_inst_U398 ( .A(aes_core_sbox_inst_n979), .Y(
        aes_core_sbox_inst_n133) );
  INVX1 aes_core_sbox_inst_U397 ( .A(aes_core_sbox_inst_n130), .Y(
        aes_core_sbox_inst_n131) );
  CLKINVX3 aes_core_sbox_inst_U396 ( .A(aes_core_sbox_inst_n2), .Y(
        aes_core_sbox_inst_n143) );
  INVX1 aes_core_sbox_inst_U395 ( .A(aes_core_sbox_inst_n602), .Y(
        aes_core_sbox_inst_n1715) );
  INVX1 aes_core_sbox_inst_U394 ( .A(aes_core_sbox_inst_n1227), .Y(
        aes_core_sbox_inst_n1597) );
  INVX1 aes_core_sbox_inst_U393 ( .A(aes_core_sbox_inst_n384), .Y(
        aes_core_sbox_inst_n141) );
  INVX1 aes_core_sbox_inst_U392 ( .A(aes_core_sbox_inst_n979), .Y(
        aes_core_sbox_inst_n132) );
  INVX1 aes_core_sbox_inst_U391 ( .A(aes_core_sbox_inst_n524), .Y(
        aes_core_sbox_inst_n1717) );
  INVX1 aes_core_sbox_inst_U390 ( .A(aes_core_sbox_inst_n1119), .Y(
        aes_core_sbox_inst_n1599) );
  INVX1 aes_core_sbox_inst_U389 ( .A(aes_core_sbox_inst_n791), .Y(
        aes_core_sbox_inst_n240) );
  CLKINVX3 aes_core_sbox_inst_U388 ( .A(aes_core_sbox_inst_n1), .Y(
        aes_core_sbox_inst_n134) );
  CLKBUFX16 aes_core_sbox_inst_U387 ( .A(aes_core_n4), .Y(
        aes_core_sbox_inst_n55) );
  AND2X1 aes_core_sbox_inst_U386 ( .A(aes_core_sbox_inst_n344), .B(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n369) );
  NOR2X2 aes_core_sbox_inst_U385 ( .A(aes_core_sbox_inst_n35), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n10) );
  INVX4 aes_core_sbox_inst_U384 ( .A(aes_core_n29), .Y(aes_core_sbox_inst_n251) );
  BUFX12 aes_core_sbox_inst_U383 ( .A(aes_core_sbox_inst_n667), .Y(
        aes_core_sbox_inst_n116) );
  BUFX1 aes_core_sbox_inst_U382 ( .A(aes_core_sbox_inst_n1679), .Y(
        aes_core_sbox_inst_n47) );
  AND2X1 aes_core_sbox_inst_U381 ( .A(aes_core_sbox_inst_n828), .B(
        aes_core_sbox_inst_n160), .Y(aes_core_sbox_inst_n890) );
  AND2X1 aes_core_sbox_inst_U380 ( .A(aes_core_sbox_inst_n1156), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1248) );
  BUFX1 aes_core_sbox_inst_U379 ( .A(aes_core_sbox_inst_n1614), .Y(
        aes_core_sbox_inst_n27) );
  BUFX1 aes_core_sbox_inst_U378 ( .A(aes_core_sbox_inst_n1676), .Y(
        aes_core_sbox_inst_n43) );
  BUFX2 aes_core_sbox_inst_U377 ( .A(aes_core_sbox_inst_n1674), .Y(
        aes_core_sbox_inst_n39) );
  INVX8 aes_core_sbox_inst_U376 ( .A(aes_core_sbox_inst_n92), .Y(
        aes_core_sbox_inst_n1585) );
  AND3X1 aes_core_sbox_inst_U375 ( .A(aes_core_sbox_inst_n310), .B(
        aes_core_sbox_inst_n311), .C(aes_core_sbox_inst_n312), .Y(
        aes_core_sbox_inst_n309) );
  BUFX12 aes_core_sbox_inst_U374 ( .A(aes_core_sbox_inst_n402), .Y(
        aes_core_sbox_inst_n65) );
  INVX8 aes_core_sbox_inst_U373 ( .A(aes_core_sbox_inst_n111), .Y(
        aes_core_sbox_inst_n248) );
  CLKBUFX2 aes_core_sbox_inst_U372 ( .A(aes_core_sbox_inst_n1675), .Y(
        aes_core_sbox_inst_n41) );
  NOR2X2 aes_core_sbox_inst_U371 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n187), .Y(aes_core_sbox_inst_n399) );
  NOR2X4 aes_core_sbox_inst_U370 ( .A(aes_core_sbox_inst_n51), .B(
        aes_core_sbox_inst_n1712), .Y(aes_core_sbox_inst_n409) );
  NOR2X4 aes_core_sbox_inst_U369 ( .A(aes_core_sbox_inst_n18), .B(
        aes_core_sbox_inst_n235), .Y(aes_core_sbox_inst_n642) );
  NOR2X1 aes_core_sbox_inst_U368 ( .A(aes_core_sbox_inst_n163), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n8) );
  NOR2X1 aes_core_sbox_inst_U367 ( .A(aes_core_sbox_inst_n177), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n7) );
  NOR2X1 aes_core_sbox_inst_U366 ( .A(aes_core_sbox_inst_n202), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n6) );
  NOR2X1 aes_core_sbox_inst_U365 ( .A(aes_core_sbox_inst_n202), .B(
        aes_core_sbox_inst_n191), .Y(aes_core_sbox_inst_n5) );
  NOR2X1 aes_core_sbox_inst_U364 ( .A(aes_core_sbox_inst_n177), .B(
        aes_core_sbox_inst_n169), .Y(aes_core_sbox_inst_n4) );
  AND2X1 aes_core_sbox_inst_U363 ( .A(aes_core_sbox_inst_n870), .B(
        aes_core_sbox_inst_n117), .Y(aes_core_sbox_inst_n697) );
  AND2X1 aes_core_sbox_inst_U362 ( .A(aes_core_sbox_inst_n1228), .B(
        aes_core_sbox_inst_n121), .Y(aes_core_sbox_inst_n1059) );
  AND2X1 aes_core_sbox_inst_U361 ( .A(aes_core_sbox_inst_n603), .B(
        aes_core_sbox_inst_n126), .Y(aes_core_sbox_inst_n464) );
  INVX8 aes_core_sbox_inst_U360 ( .A(aes_core_sbox_inst_n113), .Y(
        aes_core_sbox_inst_n225) );
  INVX8 aes_core_sbox_inst_U359 ( .A(aes_core_sbox_inst_n75), .Y(
        aes_core_sbox_inst_n1702) );
  NOR2X4 aes_core_sbox_inst_U358 ( .A(aes_core_sbox_inst_n134), .B(
        aes_core_sbox_inst_n670), .Y(aes_core_sbox_inst_n619) );
  BUFX16 aes_core_sbox_inst_U357 ( .A(aes_core_sbox_inst_n619), .Y(
        aes_core_sbox_inst_n109) );
  CLKINVX2 aes_core_sbox_inst_U356 ( .A(aes_core_sbox_inst_n69), .Y(
        aes_core_sbox_inst_n127) );
  CLKINVX2 aes_core_sbox_inst_U355 ( .A(aes_core_sbox_inst_n95), .Y(
        aes_core_sbox_inst_n122) );
  CLKBUFX2 aes_core_sbox_inst_U354 ( .A(aes_core_sbox_inst_n1616), .Y(
        aes_core_sbox_inst_n29) );
  CLKBUFX2 aes_core_sbox_inst_U353 ( .A(aes_core_sbox_inst_n1734), .Y(
        aes_core_sbox_inst_n53) );
  BUFX3 aes_core_sbox_inst_U352 ( .A(aes_core_n20), .Y(aes_core_sbox_inst_n60)
         );
  CLKBUFX16 aes_core_sbox_inst_U351 ( .A(aes_core_n22), .Y(
        aes_core_sbox_inst_n61) );
  INVX1 aes_core_sbox_inst_U350 ( .A(aes_core_n17), .Y(
        aes_core_sbox_inst_n1620) );
  NOR2X1 aes_core_sbox_inst_U349 ( .A(aes_core_sbox_inst_n180), .B(
        aes_core_n16), .Y(aes_core_sbox_inst_n1374) );
  INVX1 aes_core_sbox_inst_U348 ( .A(aes_core_n16), .Y(
        aes_core_sbox_inst_n1623) );
  INVX1 aes_core_sbox_inst_U347 ( .A(aes_core_n9), .Y(aes_core_sbox_inst_n1682) );
  INVX1 aes_core_sbox_inst_U346 ( .A(aes_core_n33), .Y(aes_core_sbox_inst_n206) );
  NOR2X1 aes_core_sbox_inst_U345 ( .A(aes_core_sbox_inst_n189), .B(
        aes_core_sbox_inst_n56), .Y(aes_core_sbox_inst_n440) );
  INVX1 aes_core_sbox_inst_U344 ( .A(aes_core_n25), .Y(aes_core_sbox_inst_n450) );
  NOR2X1 aes_core_sbox_inst_U343 ( .A(aes_core_sbox_inst_n1674), .B(
        aes_core_n13), .Y(aes_core_sbox_inst_n344) );
  NOR2X1 aes_core_sbox_inst_U342 ( .A(aes_core_sbox_inst_n36), .B(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n1455) );
  INVX1 aes_core_sbox_inst_U341 ( .A(aes_core_sbox_inst_n64), .Y(
        aes_core_sbox_inst_n209) );
  INVX1 aes_core_sbox_inst_U340 ( .A(aes_core_sbox_inst_n62), .Y(
        aes_core_sbox_inst_n1567) );
  INVX1 aes_core_sbox_inst_U339 ( .A(aes_core_sbox_inst_n56), .Y(
        aes_core_sbox_inst_n1685) );
  NAND4X1 aes_core_sbox_inst_U338 ( .A(aes_core_sbox_inst_n553), .B(
        aes_core_sbox_inst_n395), .C(aes_core_sbox_inst_n554), .D(
        aes_core_sbox_inst_n555), .Y(aes_core_sbox_inst_n552) );
  OAI2BB1X1 aes_core_sbox_inst_U337 ( .A0N(aes_core_sbox_inst_n58), .A1N(
        aes_core_sbox_inst_n89), .B0(aes_core_sbox_inst_n1665), .Y(
        aes_core_sbox_inst_n1431) );
  AOI21X1 aes_core_sbox_inst_U336 ( .A0(aes_core_sbox_inst_n61), .A1(
        aes_core_sbox_inst_n999), .B0(aes_core_sbox_inst_n1000), .Y(
        aes_core_sbox_inst_n998) );
  AOI21X1 aes_core_sbox_inst_U335 ( .A0(aes_core_sbox_inst_n337), .A1(
        aes_core_sbox_inst_n1658), .B0(aes_core_sbox_inst_n31), .Y(
        aes_core_sbox_inst_n1438) );
  AOI31X1 aes_core_sbox_inst_U334 ( .A0(aes_core_n14), .A1(
        aes_core_sbox_inst_n1677), .A2(aes_core_sbox_inst_n1357), .B0(
        aes_core_sbox_inst_n1438), .Y(aes_core_sbox_inst_n1433) );
  NOR2X1 aes_core_sbox_inst_U333 ( .A(aes_core_sbox_inst_n189), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n488) );
  NAND4X1 aes_core_sbox_inst_U332 ( .A(aes_core_sbox_inst_n1653), .B(
        aes_core_sbox_inst_n1340), .C(aes_core_sbox_inst_n1463), .D(
        aes_core_sbox_inst_n1464), .Y(aes_core_sbox_inst_n1462) );
  AOI31X1 aes_core_sbox_inst_U331 ( .A0(aes_core_n6), .A1(
        aes_core_sbox_inst_n54), .A2(aes_core_sbox_inst_n488), .B0(
        aes_core_sbox_inst_n525), .Y(aes_core_sbox_inst_n519) );
  AOI21X1 aes_core_sbox_inst_U330 ( .A0(aes_core_sbox_inst_n1459), .A1(
        aes_core_sbox_inst_n1460), .B0(aes_core_sbox_inst_n1624), .Y(
        aes_core_sbox_inst_n1458) );
  AOI222X1 aes_core_sbox_inst_U329 ( .A0(aes_core_n16), .A1(
        aes_core_sbox_inst_n1441), .B0(aes_core_sbox_inst_n1372), .B1(
        aes_core_sbox_inst_n1442), .C0(aes_core_sbox_inst_n1374), .C1(
        aes_core_sbox_inst_n1443), .Y(aes_core_sbox_inst_n1440) );
  AOI211X1 aes_core_sbox_inst_U328 ( .A0(aes_core_n16), .A1(
        aes_core_sbox_inst_n1457), .B0(aes_core_sbox_inst_n1626), .C0(
        aes_core_sbox_inst_n1458), .Y(aes_core_sbox_inst_n1439) );
  OAI22X1 aes_core_sbox_inst_U327 ( .A0(aes_core_n17), .A1(
        aes_core_sbox_inst_n1439), .B0(aes_core_sbox_inst_n1440), .B1(
        aes_core_sbox_inst_n1620), .Y(aes_core_new_sboxw[12]) );
  AOI31X1 aes_core_sbox_inst_U326 ( .A0(aes_core_sbox_inst_n1194), .A1(
        aes_core_sbox_inst_n1195), .A2(aes_core_sbox_inst_n1196), .B0(
        aes_core_sbox_inst_n316), .Y(aes_core_sbox_inst_n1193) );
  AOI21X1 aes_core_sbox_inst_U325 ( .A0(aes_core_sbox_inst_n1207), .A1(
        aes_core_sbox_inst_n1208), .B0(aes_core_n25), .Y(
        aes_core_sbox_inst_n1192) );
  AOI211X1 aes_core_sbox_inst_U324 ( .A0(aes_core_sbox_inst_n1190), .A1(
        aes_core_sbox_inst_n1191), .B0(aes_core_sbox_inst_n1192), .C0(
        aes_core_sbox_inst_n1193), .Y(aes_core_sbox_inst_n1189) );
  INVX1 aes_core_sbox_inst_U323 ( .A(aes_core_sbox_inst_n1189), .Y(
        aes_core_new_sboxw[19]) );
  AOI31X1 aes_core_sbox_inst_U322 ( .A0(aes_core_sbox_inst_n569), .A1(
        aes_core_sbox_inst_n570), .A2(aes_core_sbox_inst_n571), .B0(
        aes_core_sbox_inst_n1681), .Y(aes_core_sbox_inst_n568) );
  AOI21X1 aes_core_sbox_inst_U321 ( .A0(aes_core_sbox_inst_n582), .A1(
        aes_core_sbox_inst_n583), .B0(aes_core_n9), .Y(aes_core_sbox_inst_n567) );
  AOI211X1 aes_core_sbox_inst_U320 ( .A0(aes_core_sbox_inst_n565), .A1(
        aes_core_sbox_inst_n566), .B0(aes_core_sbox_inst_n567), .C0(
        aes_core_sbox_inst_n568), .Y(aes_core_sbox_inst_n564) );
  INVX1 aes_core_sbox_inst_U319 ( .A(aes_core_sbox_inst_n564), .Y(
        aes_core_new_sboxw[3]) );
  AOI21X1 aes_core_sbox_inst_U318 ( .A0(aes_core_sbox_inst_n849), .A1(
        aes_core_sbox_inst_n850), .B0(aes_core_n33), .Y(
        aes_core_sbox_inst_n834) );
  AOI31X1 aes_core_sbox_inst_U317 ( .A0(aes_core_sbox_inst_n1475), .A1(
        aes_core_sbox_inst_n1476), .A2(aes_core_sbox_inst_n1477), .B0(
        aes_core_sbox_inst_n1619), .Y(aes_core_sbox_inst_n1474) );
  AOI211X1 aes_core_sbox_inst_U316 ( .A0(aes_core_sbox_inst_n292), .A1(
        aes_core_sbox_inst_n125), .B0(aes_core_sbox_inst_n1479), .C0(
        aes_core_sbox_inst_n1480), .Y(aes_core_sbox_inst_n1477) );
  AOI21X1 aes_core_sbox_inst_U315 ( .A0(aes_core_sbox_inst_n404), .A1(
        aes_core_sbox_inst_n512), .B0(aes_core_sbox_inst_n423), .Y(
        aes_core_sbox_inst_n503) );
  NAND4X1 aes_core_sbox_inst_U314 ( .A(aes_core_sbox_inst_n1715), .B(
        aes_core_sbox_inst_n502), .C(aes_core_sbox_inst_n503), .D(
        aes_core_sbox_inst_n504), .Y(aes_core_sbox_inst_n501) );
  AOI211X1 aes_core_sbox_inst_U313 ( .A0(aes_core_sbox_inst_n76), .A1(
        aes_core_sbox_inst_n126), .B0(aes_core_sbox_inst_n505), .C0(
        aes_core_sbox_inst_n506), .Y(aes_core_sbox_inst_n504) );
  NOR2X1 aes_core_sbox_inst_U312 ( .A(aes_core_sbox_inst_n168), .B(
        aes_core_sbox_inst_n60), .Y(aes_core_sbox_inst_n1083) );
  NOR4BX1 aes_core_sbox_inst_U311 ( .AN(aes_core_sbox_inst_n1349), .B(
        aes_core_sbox_inst_n1350), .C(aes_core_sbox_inst_n1351), .D(
        aes_core_sbox_inst_n1352), .Y(aes_core_sbox_inst_n1325) );
  AOI211X1 aes_core_sbox_inst_U310 ( .A0(aes_core_sbox_inst_n263), .A1(
        aes_core_sbox_inst_n1327), .B0(aes_core_sbox_inst_n1328), .C0(
        aes_core_sbox_inst_n1329), .Y(aes_core_sbox_inst_n1326) );
  NOR3BX1 aes_core_sbox_inst_U309 ( .AN(aes_core_sbox_inst_n1359), .B(
        aes_core_sbox_inst_n1360), .C(aes_core_sbox_inst_n1361), .Y(
        aes_core_sbox_inst_n1324) );
  OAI222X1 aes_core_sbox_inst_U308 ( .A0(aes_core_sbox_inst_n1324), .A1(
        aes_core_sbox_inst_n1618), .B0(aes_core_sbox_inst_n1325), .B1(
        aes_core_sbox_inst_n1619), .C0(aes_core_n17), .C1(
        aes_core_sbox_inst_n1326), .Y(aes_core_new_sboxw[15]) );
  NOR4BX1 aes_core_sbox_inst_U307 ( .AN(aes_core_sbox_inst_n412), .B(
        aes_core_sbox_inst_n413), .C(aes_core_sbox_inst_n414), .D(
        aes_core_sbox_inst_n415), .Y(aes_core_sbox_inst_n372) );
  AOI211X1 aes_core_sbox_inst_U306 ( .A0(aes_core_sbox_inst_n374), .A1(
        aes_core_sbox_inst_n375), .B0(aes_core_sbox_inst_n376), .C0(
        aes_core_sbox_inst_n377), .Y(aes_core_sbox_inst_n373) );
  NOR3BX1 aes_core_sbox_inst_U305 ( .AN(aes_core_sbox_inst_n426), .B(
        aes_core_sbox_inst_n427), .C(aes_core_sbox_inst_n428), .Y(
        aes_core_sbox_inst_n371) );
  OAI222X1 aes_core_sbox_inst_U304 ( .A0(aes_core_sbox_inst_n371), .A1(
        aes_core_sbox_inst_n1680), .B0(aes_core_sbox_inst_n372), .B1(
        aes_core_sbox_inst_n1681), .C0(aes_core_n9), .C1(
        aes_core_sbox_inst_n373), .Y(aes_core_new_sboxw[7]) );
  NOR3BX1 aes_core_sbox_inst_U303 ( .AN(aes_core_sbox_inst_n1021), .B(
        aes_core_sbox_inst_n1022), .C(aes_core_sbox_inst_n1023), .Y(
        aes_core_sbox_inst_n966) );
  OAI222X1 aes_core_sbox_inst_U302 ( .A0(aes_core_sbox_inst_n966), .A1(
        aes_core_sbox_inst_n273), .B0(aes_core_sbox_inst_n967), .B1(
        aes_core_sbox_inst_n316), .C0(aes_core_n25), .C1(
        aes_core_sbox_inst_n968), .Y(aes_core_new_sboxw[23]) );
  NOR4BX1 aes_core_sbox_inst_U301 ( .AN(aes_core_sbox_inst_n1007), .B(
        aes_core_sbox_inst_n1008), .C(aes_core_sbox_inst_n1009), .D(
        aes_core_sbox_inst_n1010), .Y(aes_core_sbox_inst_n967) );
  AOI21X1 aes_core_sbox_inst_U300 ( .A0(aes_core_sbox_inst_n816), .A1(
        aes_core_sbox_inst_n817), .B0(aes_core_sbox_inst_n210), .Y(
        aes_core_sbox_inst_n815) );
  AOI222X1 aes_core_sbox_inst_U299 ( .A0(aes_core_sbox_inst_n184), .A1(
        aes_core_sbox_inst_n363), .B0(aes_core_sbox_inst_n364), .B1(
        aes_core_sbox_inst_n181), .C0(aes_core_sbox_inst_n352), .C1(
        aes_core_sbox_inst_n43), .Y(aes_core_sbox_inst_n362) );
  OAI211X1 aes_core_sbox_inst_U298 ( .A0(aes_core_sbox_inst_n47), .A1(
        aes_core_sbox_inst_n338), .B0(aes_core_sbox_inst_n361), .C0(
        aes_core_sbox_inst_n362), .Y(aes_core_sbox_inst_n347) );
  INVX1 aes_core_sbox_inst_U297 ( .A(aes_core_sbox_inst_n370), .Y(
        aes_core_sbox_inst_n1634) );
  AOI31X1 aes_core_sbox_inst_U296 ( .A0(aes_core_sbox_inst_n61), .A1(
        aes_core_sbox_inst_n30), .A2(aes_core_sbox_inst_n1083), .B0(
        aes_core_sbox_inst_n1120), .Y(aes_core_sbox_inst_n1114) );
  AOI21X1 aes_core_sbox_inst_U295 ( .A0(aes_core_sbox_inst_n549), .A1(
        aes_core_sbox_inst_n550), .B0(aes_core_sbox_inst_n1686), .Y(
        aes_core_sbox_inst_n548) );
  AOI222X1 aes_core_sbox_inst_U294 ( .A0(aes_core_sbox_inst_n56), .A1(
        aes_core_sbox_inst_n528), .B0(aes_core_sbox_inst_n529), .B1(
        aes_core_sbox_inst_n530), .C0(aes_core_sbox_inst_n440), .C1(
        aes_core_sbox_inst_n531), .Y(aes_core_sbox_inst_n527) );
  AOI211X1 aes_core_sbox_inst_U293 ( .A0(aes_core_sbox_inst_n56), .A1(
        aes_core_sbox_inst_n547), .B0(aes_core_sbox_inst_n1688), .C0(
        aes_core_sbox_inst_n548), .Y(aes_core_sbox_inst_n526) );
  OAI22X1 aes_core_sbox_inst_U292 ( .A0(aes_core_n9), .A1(
        aes_core_sbox_inst_n526), .B0(aes_core_sbox_inst_n527), .B1(
        aes_core_sbox_inst_n1682), .Y(aes_core_new_sboxw[4]) );
  AOI21X1 aes_core_sbox_inst_U291 ( .A0(aes_core_sbox_inst_n1144), .A1(
        aes_core_sbox_inst_n1145), .B0(aes_core_sbox_inst_n1568), .Y(
        aes_core_sbox_inst_n1143) );
  AOI222X1 aes_core_sbox_inst_U290 ( .A0(aes_core_sbox_inst_n62), .A1(
        aes_core_sbox_inst_n1123), .B0(aes_core_sbox_inst_n1124), .B1(
        aes_core_sbox_inst_n1125), .C0(aes_core_sbox_inst_n1035), .C1(
        aes_core_sbox_inst_n1126), .Y(aes_core_sbox_inst_n1122) );
  AOI211X1 aes_core_sbox_inst_U289 ( .A0(aes_core_sbox_inst_n62), .A1(
        aes_core_sbox_inst_n1142), .B0(aes_core_sbox_inst_n1570), .C0(
        aes_core_sbox_inst_n1143), .Y(aes_core_sbox_inst_n1121) );
  OAI22X1 aes_core_sbox_inst_U288 ( .A0(aes_core_n25), .A1(
        aes_core_sbox_inst_n1121), .B0(aes_core_sbox_inst_n1122), .B1(
        aes_core_sbox_inst_n450), .Y(aes_core_new_sboxw[20]) );
  NAND4X1 aes_core_sbox_inst_U287 ( .A(aes_core_sbox_inst_n284), .B(
        aes_core_sbox_inst_n285), .C(aes_core_sbox_inst_n286), .D(
        aes_core_sbox_inst_n287), .Y(aes_core_sbox_inst_n262) );
  AOI211X1 aes_core_sbox_inst_U286 ( .A0(aes_core_sbox_inst_n297), .A1(
        aes_core_sbox_inst_n1623), .B0(aes_core_sbox_inst_n298), .C0(
        aes_core_sbox_inst_n299), .Y(aes_core_sbox_inst_n260) );
  AOI222X1 aes_core_sbox_inst_U285 ( .A0(aes_core_sbox_inst_n262), .A1(
        aes_core_sbox_inst_n1623), .B0(aes_core_sbox_inst_n263), .B1(
        aes_core_sbox_inst_n264), .C0(aes_core_sbox_inst_n265), .C1(
        aes_core_sbox_inst_n266), .Y(aes_core_sbox_inst_n261) );
  OAI22X1 aes_core_sbox_inst_U284 ( .A0(aes_core_sbox_inst_n260), .A1(
        aes_core_sbox_inst_n1620), .B0(aes_core_n17), .B1(
        aes_core_sbox_inst_n261), .Y(aes_core_new_sboxw[9]) );
  OAI222X1 aes_core_sbox_inst_U283 ( .A0(aes_core_sbox_inst_n325), .A1(
        aes_core_sbox_inst_n1623), .B0(aes_core_sbox_inst_n1646), .B1(
        aes_core_sbox_inst_n1622), .C0(aes_core_n16), .C1(
        aes_core_sbox_inst_n326), .Y(aes_core_sbox_inst_n324) );
  OAI2BB2X1 aes_core_sbox_inst_U282 ( .B0(aes_core_n17), .B1(
        aes_core_sbox_inst_n323), .A0N(aes_core_n17), .A1N(
        aes_core_sbox_inst_n324), .Y(aes_core_new_sboxw[8]) );
  INVX1 aes_core_sbox_inst_U281 ( .A(aes_core_sbox_inst_n335), .Y(
        aes_core_sbox_inst_n1646) );
  BUFX16 aes_core_sbox_inst_U280 ( .A(aes_core_sbox_inst_n251), .Y(
        aes_core_sbox_inst_n17) );
  INVX1 aes_core_sbox_inst_U279 ( .A(aes_core_sbox_inst_n182), .Y(
        aes_core_sbox_inst_n184) );
  NOR2X1 aes_core_sbox_inst_U278 ( .A(aes_core_sbox_inst_n1620), .B(
        aes_core_sbox_inst_n1623), .Y(aes_core_sbox_inst_n1471) );
  INVX1 aes_core_sbox_inst_U277 ( .A(aes_core_sbox_inst_n1478), .Y(
        aes_core_sbox_inst_n1619) );
  INVX1 aes_core_sbox_inst_U276 ( .A(aes_core_sbox_inst_n572), .Y(
        aes_core_sbox_inst_n1681) );
  INVX1 aes_core_sbox_inst_U275 ( .A(aes_core_sbox_inst_n839), .Y(
        aes_core_sbox_inst_n205) );
  NAND2BX1 aes_core_sbox_inst_U274 ( .AN(aes_core_sbox_inst_n368), .B(
        aes_core_sbox_inst_n45), .Y(aes_core_sbox_inst_n1395) );
  INVX1 aes_core_sbox_inst_U273 ( .A(aes_core_sbox_inst_n1197), .Y(
        aes_core_sbox_inst_n316) );
  NAND2X1 aes_core_sbox_inst_U272 ( .A(aes_core_sbox_inst_n314), .B(
        aes_core_sbox_inst_n80), .Y(aes_core_sbox_inst_n1412) );
  NOR2X1 aes_core_sbox_inst_U271 ( .A(aes_core_sbox_inst_n1685), .B(
        aes_core_sbox_inst_n189), .Y(aes_core_sbox_inst_n374) );
  NOR2X1 aes_core_sbox_inst_U270 ( .A(aes_core_sbox_inst_n1636), .B(
        aes_core_sbox_inst_n38), .Y(aes_core_sbox_inst_n292) );
  AND2X2 aes_core_sbox_inst_U269 ( .A(aes_core_sbox_inst_n561), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n743) );
  INVX1 aes_core_sbox_inst_U268 ( .A(aes_core_sbox_inst_n360), .Y(
        aes_core_sbox_inst_n1633) );
  NAND2X1 aes_core_sbox_inst_U267 ( .A(aes_core_sbox_inst_n1041), .B(
        aes_core_sbox_inst_n167), .Y(aes_core_sbox_inst_n1256) );
  BUFX3 aes_core_sbox_inst_U266 ( .A(aes_core_sbox_inst_n1614), .Y(
        aes_core_sbox_inst_n26) );
  INVX1 aes_core_sbox_inst_U265 ( .A(aes_core_sbox_inst_n490), .Y(
        aes_core_sbox_inst_n1730) );
  INVX1 aes_core_sbox_inst_U264 ( .A(aes_core_sbox_inst_n1085), .Y(
        aes_core_sbox_inst_n1612) );
  INVX1 aes_core_sbox_inst_U263 ( .A(aes_core_sbox_inst_n84), .Y(
        aes_core_sbox_inst_n1678) );
  INVX1 aes_core_sbox_inst_U262 ( .A(aes_core_sbox_inst_n1393), .Y(
        aes_core_sbox_inst_n1673) );
  INVX1 aes_core_sbox_inst_U261 ( .A(aes_core_sbox_inst_n796), .Y(
        aes_core_sbox_inst_n211) );
  INVX1 aes_core_sbox_inst_U260 ( .A(aes_core_sbox_inst_n529), .Y(
        aes_core_sbox_inst_n1687) );
  NOR2X1 aes_core_sbox_inst_U259 ( .A(aes_core_sbox_inst_n133), .B(
        aes_core_sbox_inst_n25), .Y(aes_core_sbox_inst_n1103) );
  NAND3X1 aes_core_sbox_inst_U258 ( .A(aes_core_sbox_inst_n471), .B(
        aes_core_sbox_inst_n189), .C(aes_core_sbox_inst_n71), .Y(
        aes_core_sbox_inst_n581) );
  NOR2X1 aes_core_sbox_inst_U257 ( .A(aes_core_sbox_inst_n1567), .B(
        aes_core_sbox_inst_n166), .Y(aes_core_sbox_inst_n969) );
  NOR2X1 aes_core_sbox_inst_U256 ( .A(aes_core_sbox_inst_n209), .B(
        aes_core_sbox_inst_n148), .Y(aes_core_sbox_inst_n607) );
  NOR2X1 aes_core_sbox_inst_U255 ( .A(aes_core_sbox_inst_n276), .B(
        aes_core_sbox_inst_n344), .Y(aes_core_sbox_inst_n1334) );
  NOR2X1 aes_core_sbox_inst_U254 ( .A(aes_core_sbox_inst_n1685), .B(
        aes_core_sbox_inst_n186), .Y(aes_core_sbox_inst_n592) );
  INVX1 aes_core_sbox_inst_U253 ( .A(aes_core_sbox_inst_n721), .Y(
        aes_core_sbox_inst_n215) );
  INVX1 aes_core_sbox_inst_U252 ( .A(aes_core_sbox_inst_n71), .Y(
        aes_core_sbox_inst_n1720) );
  NAND2X1 aes_core_sbox_inst_U251 ( .A(aes_core_sbox_inst_n446), .B(
        aes_core_sbox_inst_n188), .Y(aes_core_sbox_inst_n751) );
  INVX1 aes_core_sbox_inst_U250 ( .A(aes_core_sbox_inst_n89), .Y(
        aes_core_sbox_inst_n1664) );
  INVX1 aes_core_sbox_inst_U249 ( .A(aes_core_sbox_inst_n76), .Y(
        aes_core_sbox_inst_n1714) );
  INVX1 aes_core_sbox_inst_U248 ( .A(aes_core_sbox_inst_n90), .Y(
        aes_core_sbox_inst_n1638) );
  INVX1 aes_core_sbox_inst_U247 ( .A(aes_core_sbox_inst_n1124), .Y(
        aes_core_sbox_inst_n1569) );
  INVX1 aes_core_sbox_inst_U246 ( .A(aes_core_sbox_inst_n1205), .Y(
        aes_core_sbox_inst_n1613) );
  AOI21X1 aes_core_sbox_inst_U245 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n145), .B0(aes_core_sbox_inst_n358), .Y(
        aes_core_sbox_inst_n354) );
  INVX1 aes_core_sbox_inst_U244 ( .A(aes_core_sbox_inst_n580), .Y(
        aes_core_sbox_inst_n1731) );
  NOR2X1 aes_core_sbox_inst_U243 ( .A(aes_core_sbox_inst_n1), .B(
        aes_core_sbox_inst_n17), .Y(aes_core_sbox_inst_n775) );
  AOI221X1 aes_core_sbox_inst_U242 ( .A0(aes_core_sbox_inst_n344), .A1(
        aes_core_sbox_inst_n84), .B0(aes_core_sbox_inst_n345), .B1(
        aes_core_sbox_inst_n45), .C0(aes_core_sbox_inst_n346), .Y(
        aes_core_sbox_inst_n343) );
  NOR2X1 aes_core_sbox_inst_U241 ( .A(aes_core_sbox_inst_n561), .B(
        aes_core_sbox_inst_n538), .Y(aes_core_sbox_inst_n590) );
  NOR2X1 aes_core_sbox_inst_U240 ( .A(aes_core_sbox_inst_n1567), .B(
        aes_core_sbox_inst_n164), .Y(aes_core_sbox_inst_n1217) );
  BUFX12 aes_core_sbox_inst_U239 ( .A(aes_core_sbox_inst_n236), .Y(
        aes_core_sbox_inst_n15) );
  NAND2X1 aes_core_sbox_inst_U238 ( .A(aes_core_sbox_inst_n679), .B(
        aes_core_sbox_inst_n148), .Y(aes_core_sbox_inst_n898) );
  INVX1 aes_core_sbox_inst_U237 ( .A(aes_core_sbox_inst_n114), .Y(
        aes_core_sbox_inst_n237) );
  BUFX1 aes_core_sbox_inst_U236 ( .A(aes_core_sbox_inst_n1676), .Y(
        aes_core_sbox_inst_n42) );
  INVX1 aes_core_sbox_inst_U235 ( .A(aes_core_sbox_inst_n723), .Y(
        aes_core_sbox_inst_n253) );
  NAND4X1 aes_core_sbox_inst_U234 ( .A(aes_core_sbox_inst_n1668), .B(
        aes_core_sbox_inst_n320), .C(aes_core_sbox_inst_n1417), .D(
        aes_core_sbox_inst_n1418), .Y(aes_core_sbox_inst_n1416) );
  AOI211X1 aes_core_sbox_inst_U233 ( .A0(aes_core_sbox_inst_n89), .A1(
        aes_core_sbox_inst_n41), .B0(aes_core_sbox_inst_n1419), .C0(
        aes_core_sbox_inst_n1420), .Y(aes_core_sbox_inst_n1418) );
  INVX1 aes_core_sbox_inst_U232 ( .A(aes_core_sbox_inst_n74), .Y(
        aes_core_sbox_inst_n1706) );
  OAI211X1 aes_core_sbox_inst_U231 ( .A0(aes_core_sbox_inst_n1081), .A1(
        aes_core_sbox_inst_n1579), .B0(aes_core_sbox_inst_n1604), .C0(
        aes_core_sbox_inst_n1082), .Y(aes_core_sbox_inst_n1075) );
  INVX1 aes_core_sbox_inst_U230 ( .A(aes_core_sbox_inst_n1084), .Y(
        aes_core_sbox_inst_n1604) );
  NOR2X1 aes_core_sbox_inst_U229 ( .A(aes_core_sbox_inst_n828), .B(
        aes_core_sbox_inst_n805), .Y(aes_core_sbox_inst_n857) );
  AOI22X1 aes_core_sbox_inst_U228 ( .A0(aes_core_sbox_inst_n292), .A1(
        aes_core_sbox_inst_n42), .B0(aes_core_sbox_inst_n179), .B1(
        aes_core_sbox_inst_n1532), .Y(aes_core_sbox_inst_n1531) );
  OAI211X1 aes_core_sbox_inst_U227 ( .A0(aes_core_sbox_inst_n81), .A1(
        aes_core_sbox_inst_n1661), .B0(aes_core_sbox_inst_n1365), .C0(
        aes_core_sbox_inst_n1533), .Y(aes_core_sbox_inst_n1532) );
  INVX1 aes_core_sbox_inst_U226 ( .A(aes_core_sbox_inst_n170), .Y(
        aes_core_sbox_inst_n171) );
  INVX1 aes_core_sbox_inst_U225 ( .A(aes_core_sbox_inst_n174), .Y(
        aes_core_sbox_inst_n175) );
  NOR2X1 aes_core_sbox_inst_U224 ( .A(aes_core_sbox_inst_n1623), .B(
        aes_core_sbox_inst_n180), .Y(aes_core_sbox_inst_n263) );
  INVX1 aes_core_sbox_inst_U223 ( .A(aes_core_sbox_inst_n1484), .Y(
        aes_core_sbox_inst_n1627) );
  INVX1 aes_core_sbox_inst_U222 ( .A(aes_core_sbox_inst_n565), .Y(
        aes_core_sbox_inst_n1680) );
  INVX1 aes_core_sbox_inst_U221 ( .A(aes_core_sbox_inst_n1190), .Y(
        aes_core_sbox_inst_n273) );
  INVX1 aes_core_sbox_inst_U220 ( .A(aes_core_sbox_inst_n832), .Y(
        aes_core_sbox_inst_n204) );
  INVX1 aes_core_sbox_inst_U219 ( .A(aes_core_sbox_inst_n196), .Y(
        aes_core_sbox_inst_n202) );
  BUFX3 aes_core_sbox_inst_U218 ( .A(aes_core_sbox_inst_n1677), .Y(
        aes_core_sbox_inst_n44) );
  INVX1 aes_core_sbox_inst_U217 ( .A(aes_core_sbox_inst_n508), .Y(
        aes_core_sbox_inst_n1726) );
  NOR2X1 aes_core_sbox_inst_U216 ( .A(aes_core_sbox_inst_n201), .B(
        aes_core_sbox_inst_n1703), .Y(aes_core_sbox_inst_n398) );
  INVX1 aes_core_sbox_inst_U215 ( .A(aes_core_sbox_inst_n859), .Y(
        aes_core_sbox_inst_n208) );
  INVX1 aes_core_sbox_inst_U214 ( .A(aes_core_sbox_inst_n315), .Y(
        aes_core_sbox_inst_n1637) );
  NAND3X1 aes_core_sbox_inst_U213 ( .A(aes_core_sbox_inst_n1678), .B(
        aes_core_sbox_inst_n39), .C(aes_core_sbox_inst_n1656), .Y(
        aes_core_sbox_inst_n353) );
  INVX1 aes_core_sbox_inst_U212 ( .A(aes_core_sbox_inst_n1446), .Y(
        aes_core_sbox_inst_n1656) );
  NOR2X1 aes_core_sbox_inst_U211 ( .A(aes_core_sbox_inst_n1630), .B(
        aes_core_sbox_inst_n35), .Y(aes_core_sbox_inst_n307) );
  INVX1 aes_core_sbox_inst_U210 ( .A(aes_core_n18), .Y(aes_core_sbox_inst_n177) );
  NOR2X1 aes_core_sbox_inst_U209 ( .A(aes_core_sbox_inst_n175), .B(
        aes_core_sbox_inst_n22), .Y(aes_core_sbox_inst_n993) );
  NOR2X1 aes_core_sbox_inst_U208 ( .A(aes_core_sbox_inst_n161), .B(
        aes_core_sbox_inst_n14), .Y(aes_core_sbox_inst_n631) );
  AOI21X1 aes_core_sbox_inst_U207 ( .A0(aes_core_sbox_inst_n83), .A1(
        aes_core_sbox_inst_n42), .B0(aes_core_sbox_inst_n267), .Y(
        aes_core_sbox_inst_n1403) );
  NOR2X1 aes_core_sbox_inst_U206 ( .A(aes_core_sbox_inst_n32), .B(
        aes_core_sbox_inst_n46), .Y(aes_core_sbox_inst_n1528) );
  NAND3X1 aes_core_sbox_inst_U205 ( .A(aes_core_sbox_inst_n128), .B(
        aes_core_sbox_inst_n1732), .C(aes_core_sbox_inst_n1704), .Y(
        aes_core_sbox_inst_n732) );
  NAND3X1 aes_core_sbox_inst_U204 ( .A(aes_core_sbox_inst_n123), .B(
        aes_core_sbox_inst_n27), .C(aes_core_sbox_inst_n1586), .Y(
        aes_core_sbox_inst_n1237) );
  NOR2X1 aes_core_sbox_inst_U203 ( .A(aes_core_sbox_inst_n338), .B(
        aes_core_sbox_inst_n144), .Y(aes_core_sbox_inst_n1368) );
  INVX1 aes_core_sbox_inst_U202 ( .A(aes_core_sbox_inst_n385), .Y(
        aes_core_sbox_inst_n1704) );
  NOR2X1 aes_core_sbox_inst_U201 ( .A(aes_core_sbox_inst_n1703), .B(
        aes_core_sbox_inst_n1691), .Y(aes_core_sbox_inst_n424) );
  NOR2X1 aes_core_sbox_inst_U200 ( .A(aes_core_sbox_inst_n1607), .B(
        aes_core_sbox_inst_n1573), .Y(aes_core_sbox_inst_n987) );
  NOR2X1 aes_core_sbox_inst_U199 ( .A(aes_core_sbox_inst_n1725), .B(
        aes_core_sbox_inst_n1691), .Y(aes_core_sbox_inst_n392) );
  BUFX16 aes_core_sbox_inst_U198 ( .A(aes_core_sbox_inst_n409), .Y(
        aes_core_sbox_inst_n68) );
  INVX1 aes_core_sbox_inst_U197 ( .A(aes_core_sbox_inst_n618), .Y(
        aes_core_sbox_inst_n227) );
  INVX1 aes_core_sbox_inst_U196 ( .A(aes_core_sbox_inst_n290), .Y(
        aes_core_sbox_inst_n1628) );
  INVX1 aes_core_sbox_inst_U195 ( .A(aes_core_sbox_inst_n265), .Y(
        aes_core_sbox_inst_n1622) );
  INVX1 aes_core_sbox_inst_U194 ( .A(aes_core_sbox_inst_n333), .Y(
        aes_core_sbox_inst_n1658) );
  INVX1 aes_core_sbox_inst_U193 ( .A(aes_core_sbox_inst_n1547), .Y(
        aes_core_sbox_inst_n1695) );
  INVX1 aes_core_sbox_inst_U192 ( .A(aes_core_sbox_inst_n657), .Y(
        aes_core_sbox_inst_n214) );
  INVX1 aes_core_sbox_inst_U191 ( .A(aes_core_sbox_inst_n352), .Y(
        aes_core_sbox_inst_n1632) );
  NAND2X1 aes_core_sbox_inst_U190 ( .A(aes_core_sbox_inst_n94), .B(
        aes_core_sbox_inst_n175), .Y(aes_core_sbox_inst_n990) );
  NAND2X1 aes_core_sbox_inst_U189 ( .A(aes_core_sbox_inst_n68), .B(
        aes_core_sbox_inst_n201), .Y(aes_core_sbox_inst_n395) );
  NAND2X1 aes_core_sbox_inst_U188 ( .A(aes_core_sbox_inst_n356), .B(
        aes_core_sbox_inst_n124), .Y(aes_core_sbox_inst_n320) );
  INVX1 aes_core_sbox_inst_U187 ( .A(aes_core_sbox_inst_n702), .Y(
        aes_core_sbox_inst_n222) );
  NOR2X1 aes_core_sbox_inst_U186 ( .A(aes_core_sbox_inst_n19), .B(
        aes_core_sbox_inst_n235), .Y(aes_core_sbox_inst_n843) );
  INVX1 aes_core_sbox_inst_U185 ( .A(aes_core_sbox_inst_n628), .Y(
        aes_core_sbox_inst_n234) );
  AOI21X1 aes_core_sbox_inst_U184 ( .A0(aes_core_sbox_inst_n118), .A1(
        aes_core_sbox_inst_n630), .B0(aes_core_sbox_inst_n234), .Y(
        aes_core_sbox_inst_n665) );
  NAND2X1 aes_core_sbox_inst_U183 ( .A(aes_core_sbox_inst_n108), .B(
        aes_core_sbox_inst_n163), .Y(aes_core_sbox_inst_n628) );
  INVX1 aes_core_sbox_inst_U182 ( .A(aes_core_sbox_inst_n1432), .Y(
        aes_core_sbox_inst_n1665) );
  INVX1 aes_core_sbox_inst_U181 ( .A(aes_core_sbox_inst_n1201), .Y(
        aes_core_sbox_inst_n1587) );
  INVX1 aes_core_sbox_inst_U180 ( .A(aes_core_sbox_inst_n576), .Y(
        aes_core_sbox_inst_n1705) );
  INVX1 aes_core_sbox_inst_U179 ( .A(aes_core_sbox_inst_n563), .Y(
        aes_core_sbox_inst_n1716) );
  INVX1 aes_core_sbox_inst_U178 ( .A(aes_core_sbox_inst_n470), .Y(
        aes_core_sbox_inst_n1707) );
  INVX1 aes_core_sbox_inst_U177 ( .A(aes_core_sbox_inst_n1065), .Y(
        aes_core_sbox_inst_n1589) );
  NAND4BX1 aes_core_sbox_inst_U176 ( .AN(aes_core_sbox_inst_n1139), .B(
        aes_core_sbox_inst_n989), .C(aes_core_sbox_inst_n1598), .D(
        aes_core_sbox_inst_n1130), .Y(aes_core_sbox_inst_n1137) );
  NOR2X1 aes_core_sbox_inst_U175 ( .A(aes_core_sbox_inst_n124), .B(
        aes_core_sbox_inst_n1651), .Y(aes_core_sbox_inst_n1423) );
  INVX1 aes_core_sbox_inst_U174 ( .A(aes_core_sbox_inst_n139), .Y(
        aes_core_sbox_inst_n140) );
  BUFX3 aes_core_sbox_inst_U173 ( .A(aes_core_sbox_inst_n1735), .Y(
        aes_core_sbox_inst_n54) );
  BUFX3 aes_core_sbox_inst_U172 ( .A(aes_core_sbox_inst_n1617), .Y(
        aes_core_sbox_inst_n30) );
  BUFX3 aes_core_sbox_inst_U171 ( .A(aes_core_sbox_inst_n259), .Y(
        aes_core_sbox_inst_n20) );
  NOR2X1 aes_core_sbox_inst_U170 ( .A(aes_core_sbox_inst_n121), .B(
        aes_core_sbox_inst_n1600), .Y(aes_core_sbox_inst_n1119) );
  NOR2X1 aes_core_sbox_inst_U169 ( .A(aes_core_sbox_inst_n1600), .B(
        aes_core_sbox_inst_n28), .Y(aes_core_sbox_inst_n1072) );
  CLKINVX3 aes_core_sbox_inst_U168 ( .A(aes_core_sbox_inst_n120), .Y(
        aes_core_sbox_inst_n118) );
  BUFX3 aes_core_sbox_inst_U167 ( .A(aes_core_sbox_inst_n1616), .Y(
        aes_core_sbox_inst_n28) );
  INVX1 aes_core_sbox_inst_U166 ( .A(aes_core_sbox_inst_n869), .Y(
        aes_core_sbox_inst_n238) );
  CLKINVX3 aes_core_sbox_inst_U165 ( .A(aes_core_sbox_inst_n137), .Y(
        aes_core_sbox_inst_n139) );
  CLKINVX3 aes_core_sbox_inst_U164 ( .A(aes_core_sbox_inst_n133), .Y(
        aes_core_sbox_inst_n130) );
  CLKINVX3 aes_core_sbox_inst_U163 ( .A(aes_core_sbox_inst_n1), .Y(
        aes_core_sbox_inst_n135) );
  BUFX12 aes_core_sbox_inst_U162 ( .A(aes_core_sbox_inst_n434), .Y(
        aes_core_sbox_inst_n78) );
  AOI31X2 aes_core_sbox_inst_U161 ( .A0(aes_core_sbox_inst_n836), .A1(
        aes_core_sbox_inst_n837), .A2(aes_core_sbox_inst_n838), .B0(
        aes_core_sbox_inst_n205), .Y(aes_core_sbox_inst_n835) );
  NOR2X4 aes_core_sbox_inst_U160 ( .A(aes_core_sbox_inst_n46), .B(
        aes_core_sbox_inst_n58), .Y(aes_core_sbox_inst_n327) );
  INVX4 aes_core_sbox_inst_U159 ( .A(aes_core_n13), .Y(
        aes_core_sbox_inst_n1672) );
  INVX4 aes_core_sbox_inst_U158 ( .A(aes_core_n21), .Y(
        aes_core_sbox_inst_n1610) );
  INVX1 aes_core_sbox_inst_U157 ( .A(aes_core_sbox_inst_n847), .Y(
        aes_core_sbox_inst_n254) );
  NOR2X4 aes_core_sbox_inst_U156 ( .A(aes_core_sbox_inst_n145), .B(
        aes_core_sbox_inst_n38), .Y(aes_core_sbox_inst_n313) );
  NOR2X1 aes_core_sbox_inst_U155 ( .A(aes_core_sbox_inst_n221), .B(
        aes_core_sbox_inst_n17), .Y(aes_core_sbox_inst_n840) );
  INVX8 aes_core_sbox_inst_U154 ( .A(aes_core_sbox_inst_n73), .Y(
        aes_core_sbox_inst_n1725) );
  INVX8 aes_core_sbox_inst_U153 ( .A(aes_core_sbox_inst_n99), .Y(
        aes_core_sbox_inst_n1607) );
  NOR2X4 aes_core_sbox_inst_U152 ( .A(aes_core_sbox_inst_n243), .B(
        aes_core_sbox_inst_n18), .Y(aes_core_sbox_inst_n630) );
  BUFX2 aes_core_sbox_inst_U151 ( .A(aes_core_sbox_inst_n1675), .Y(
        aes_core_sbox_inst_n40) );
  NOR2X4 aes_core_sbox_inst_U150 ( .A(aes_core_sbox_inst_n151), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n670) );
  AOI211X2 aes_core_sbox_inst_U149 ( .A0(aes_core_sbox_inst_n614), .A1(
        aes_core_sbox_inst_n259), .B0(aes_core_sbox_inst_n654), .C0(
        aes_core_sbox_inst_n869), .Y(aes_core_sbox_inst_n868) );
  NOR2X1 aes_core_sbox_inst_U148 ( .A(aes_core_sbox_inst_n126), .B(
        aes_core_sbox_inst_n1718), .Y(aes_core_sbox_inst_n524) );
  CLKINVX3 aes_core_sbox_inst_U147 ( .A(aes_core_sbox_inst_n120), .Y(
        aes_core_sbox_inst_n119) );
  NOR2X1 aes_core_sbox_inst_U146 ( .A(aes_core_sbox_inst_n1718), .B(
        aes_core_sbox_inst_n52), .Y(aes_core_sbox_inst_n477) );
  BUFX2 aes_core_sbox_inst_U145 ( .A(aes_core_sbox_inst_n1734), .Y(
        aes_core_sbox_inst_n52) );
  BUFX16 aes_core_sbox_inst_U144 ( .A(aes_core_n11), .Y(aes_core_sbox_inst_n58) );
  NOR2X1 aes_core_sbox_inst_U143 ( .A(aes_core_sbox_inst_n182), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n1357) );
  NOR2X2 aes_core_sbox_inst_U142 ( .A(aes_core_sbox_inst_n59), .B(
        aes_core_sbox_inst_n179), .Y(aes_core_sbox_inst_n293) );
  INVX1 aes_core_sbox_inst_U141 ( .A(aes_core_sbox_inst_n102), .Y(
        aes_core_sbox_inst_n1596) );
  INVX1 aes_core_sbox_inst_U140 ( .A(aes_core_sbox_inst_n85), .Y(
        aes_core_sbox_inst_n1670) );
  NOR2X1 aes_core_sbox_inst_U139 ( .A(aes_core_sbox_inst_n1156), .B(
        aes_core_sbox_inst_n1133), .Y(aes_core_sbox_inst_n1215) );
  NOR2X1 aes_core_sbox_inst_U138 ( .A(aes_core_sbox_inst_n32), .B(
        aes_core_sbox_inst_n43), .Y(aes_core_sbox_inst_n334) );
  NOR2X1 aes_core_sbox_inst_U137 ( .A(aes_core_sbox_inst_n16), .B(
        aes_core_sbox_inst_n159), .Y(aes_core_sbox_inst_n830) );
  INVX1 aes_core_sbox_inst_U136 ( .A(aes_core_sbox_inst_n86), .Y(
        aes_core_sbox_inst_n1669) );
  BUFX3 aes_core_sbox_inst_U135 ( .A(aes_core_sbox_inst_n241), .Y(
        aes_core_sbox_inst_n16) );
  INVX1 aes_core_sbox_inst_U134 ( .A(aes_core_sbox_inst_n718), .Y(
        aes_core_sbox_inst_n231) );
  CLKINVX3 aes_core_sbox_inst_U133 ( .A(aes_core_sbox_inst_n132), .Y(
        aes_core_sbox_inst_n129) );
  CLKINVX3 aes_core_sbox_inst_U132 ( .A(aes_core_sbox_inst_n141), .Y(
        aes_core_sbox_inst_n138) );
  AOI21X1 aes_core_sbox_inst_U131 ( .A0(aes_core_n14), .A1(
        aes_core_sbox_inst_n293), .B0(aes_core_sbox_inst_n288), .Y(
        aes_core_sbox_inst_n1345) );
  BUFX3 aes_core_sbox_inst_U130 ( .A(aes_core_sbox_inst_n1610), .Y(
        aes_core_sbox_inst_n25) );
  NOR2X1 aes_core_sbox_inst_U129 ( .A(aes_core_sbox_inst_n1334), .B(
        aes_core_n14), .Y(aes_core_sbox_inst_n1380) );
  AOI22X1 aes_core_sbox_inst_U128 ( .A0(aes_core_sbox_inst_n453), .A1(
        aes_core_sbox_inst_n5), .B0(aes_core_sbox_inst_n529), .B1(
        aes_core_sbox_inst_n552), .Y(aes_core_sbox_inst_n551) );
  AOI22X1 aes_core_sbox_inst_U127 ( .A0(aes_core_sbox_inst_n291), .A1(
        aes_core_sbox_inst_n80), .B0(aes_core_sbox_inst_n1372), .B1(
        aes_core_sbox_inst_n1462), .Y(aes_core_sbox_inst_n1461) );
  INVX1 aes_core_sbox_inst_U126 ( .A(aes_core_sbox_inst_n97), .Y(
        aes_core_sbox_inst_n1602) );
  BUFX3 aes_core_sbox_inst_U125 ( .A(aes_core_sbox_inst_n1602), .Y(
        aes_core_sbox_inst_n24) );
  INVX1 aes_core_sbox_inst_U124 ( .A(aes_core_sbox_inst_n980), .Y(
        aes_core_sbox_inst_n1586) );
  INVX1 aes_core_sbox_inst_U123 ( .A(aes_core_sbox_inst_n1429), .Y(
        aes_core_sbox_inst_n1631) );
  NAND3X1 aes_core_sbox_inst_U122 ( .A(aes_core_sbox_inst_n119), .B(
        aes_core_sbox_inst_n18), .C(aes_core_sbox_inst_n227), .Y(
        aes_core_sbox_inst_n879) );
  NOR2X1 aes_core_sbox_inst_U121 ( .A(aes_core_sbox_inst_n40), .B(
        aes_core_sbox_inst_n1660), .Y(aes_core_sbox_inst_n1398) );
  NOR2X1 aes_core_sbox_inst_U120 ( .A(aes_core_sbox_inst_n1723), .B(
        aes_core_sbox_inst_n126), .Y(aes_core_sbox_inst_n489) );
  NOR2X1 aes_core_sbox_inst_U119 ( .A(aes_core_sbox_inst_n1605), .B(
        aes_core_sbox_inst_n121), .Y(aes_core_sbox_inst_n1084) );
  NOR2X1 aes_core_sbox_inst_U118 ( .A(aes_core_sbox_inst_n246), .B(
        aes_core_sbox_inst_n117), .Y(aes_core_sbox_inst_n722) );
  NOR2X1 aes_core_sbox_inst_U117 ( .A(aes_core_sbox_inst_n1600), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1158) );
  INVX1 aes_core_sbox_inst_U116 ( .A(aes_core_sbox_inst_n1064), .Y(
        aes_core_sbox_inst_n1580) );
  NOR2X1 aes_core_sbox_inst_U115 ( .A(aes_core_sbox_inst_n36), .B(
        aes_core_sbox_inst_n143), .Y(aes_core_sbox_inst_n1425) );
  NOR2X1 aes_core_sbox_inst_U114 ( .A(aes_core_sbox_inst_n32), .B(
        aes_core_sbox_inst_n124), .Y(aes_core_sbox_inst_n267) );
  INVX1 aes_core_sbox_inst_U113 ( .A(aes_core_sbox_inst_n437), .Y(
        aes_core_sbox_inst_n128) );
  INVX1 aes_core_sbox_inst_U112 ( .A(aes_core_sbox_inst_n1032), .Y(
        aes_core_sbox_inst_n123) );
  INVX1 aes_core_sbox_inst_U111 ( .A(aes_core_sbox_inst_n1461), .Y(
        aes_core_sbox_inst_n1626) );
  BUFX4 aes_core_sbox_inst_U110 ( .A(aes_core_sbox_inst_n1663), .Y(
        aes_core_sbox_inst_n35) );
  INVX1 aes_core_sbox_inst_U109 ( .A(aes_core_sbox_inst_n100), .Y(
        aes_core_sbox_inst_n1588) );
  NOR2X1 aes_core_sbox_inst_U108 ( .A(aes_core_sbox_inst_n39), .B(
        aes_core_sbox_inst_n179), .Y(aes_core_sbox_inst_n359) );
  INVX1 aes_core_sbox_inst_U107 ( .A(aes_core_sbox_inst_n1305), .Y(
        aes_core_sbox_inst_n1577) );
  NOR2X2 aes_core_sbox_inst_U106 ( .A(aes_core_sbox_inst_n1215), .B(
        aes_core_sbox_inst_n61), .Y(aes_core_sbox_inst_n1041) );
  BUFX3 aes_core_sbox_inst_U105 ( .A(aes_core_sbox_inst_n1679), .Y(
        aes_core_sbox_inst_n46) );
  NOR2X4 aes_core_sbox_inst_U104 ( .A(aes_core_sbox_inst_n1645), .B(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n356) );
  NOR2X4 aes_core_sbox_inst_U103 ( .A(aes_core_sbox_inst_n129), .B(
        aes_core_sbox_inst_n95), .Y(aes_core_sbox_inst_n981) );
  BUFX3 aes_core_sbox_inst_U102 ( .A(aes_core_sbox_inst_n1669), .Y(
        aes_core_sbox_inst_n36) );
  CLKBUFX8 aes_core_sbox_inst_U101 ( .A(aes_core_sbox_inst_n327), .Y(
        aes_core_sbox_inst_n80) );
  NOR2X1 aes_core_sbox_inst_U100 ( .A(aes_core_sbox_inst_n63), .B(
        aes_core_sbox_inst_n146), .Y(aes_core_sbox_inst_n637) );
  NOR2X4 aes_core_sbox_inst_U99 ( .A(aes_core_sbox_inst_n34), .B(aes_core_n13), 
        .Y(aes_core_sbox_inst_n321) );
  NOR2X2 aes_core_sbox_inst_U98 ( .A(aes_core_sbox_inst_n33), .B(
        aes_core_sbox_inst_n59), .Y(aes_core_sbox_inst_n272) );
  BUFX3 aes_core_sbox_inst_U97 ( .A(aes_core_sbox_inst_n1732), .Y(
        aes_core_sbox_inst_n51) );
  BUFX12 aes_core_sbox_inst_U96 ( .A(aes_core_sbox_inst_n305), .Y(
        aes_core_sbox_inst_n87) );
  CLKINVX1 aes_core_sbox_inst_U95 ( .A(aes_core_n19), .Y(
        aes_core_sbox_inst_n172) );
  INVX4 aes_core_sbox_inst_U94 ( .A(aes_core_sbox_inst_n203), .Y(
        aes_core_sbox_inst_n199) );
  NOR2X4 aes_core_sbox_inst_U93 ( .A(aes_core_sbox_inst_n33), .B(
        aes_core_sbox_inst_n39), .Y(aes_core_sbox_inst_n274) );
  NOR2X2 aes_core_sbox_inst_U92 ( .A(aes_core_sbox_inst_n117), .B(
        aes_core_sbox_inst_n232), .Y(aes_core_sbox_inst_n654) );
  BUFX3 aes_core_sbox_inst_U91 ( .A(aes_core_sbox_inst_n437), .Y(
        aes_core_sbox_inst_n69) );
  BUFX3 aes_core_sbox_inst_U90 ( .A(aes_core_sbox_inst_n1032), .Y(
        aes_core_sbox_inst_n95) );
  NOR2X2 aes_core_sbox_inst_U89 ( .A(aes_core_sbox_inst_n169), .B(
        aes_core_sbox_inst_n174), .Y(aes_core_sbox_inst_n1032) );
  CLKINVX3 aes_core_sbox_inst_U88 ( .A(aes_core_sbox_inst_n63), .Y(
        aes_core_sbox_inst_n255) );
  INVX2 aes_core_sbox_inst_U87 ( .A(aes_core_sbox_inst_n98), .Y(
        aes_core_sbox_inst_n1600) );
  NOR2X1 aes_core_sbox_inst_U86 ( .A(aes_core_sbox_inst_n176), .B(
        aes_core_sbox_inst_n173), .Y(aes_core_sbox_inst_n979) );
  INVX1 aes_core_sbox_inst_U85 ( .A(aes_core_n18), .Y(aes_core_sbox_inst_n176)
         );
  NOR2X2 aes_core_sbox_inst_U84 ( .A(aes_core_sbox_inst_n1703), .B(
        aes_core_sbox_inst_n55), .Y(aes_core_sbox_inst_n3) );
  CLKINVX3 aes_core_sbox_inst_U83 ( .A(aes_core_sbox_inst_n158), .Y(
        aes_core_sbox_inst_n159) );
  BUFX3 aes_core_sbox_inst_U82 ( .A(aes_core_sbox_inst_n257), .Y(
        aes_core_sbox_inst_n19) );
  INVX1 aes_core_sbox_inst_U81 ( .A(aes_core_sbox_inst_n157), .Y(
        aes_core_sbox_inst_n163) );
  INVX1 aes_core_sbox_inst_U80 ( .A(aes_core_n2), .Y(aes_core_sbox_inst_n198)
         );
  INVX1 aes_core_sbox_inst_U79 ( .A(aes_core_n26), .Y(aes_core_sbox_inst_n158)
         );
  INVX1 aes_core_sbox_inst_U78 ( .A(aes_core_n31), .Y(aes_core_sbox_inst_n150)
         );
  CLKINVX3 aes_core_sbox_inst_U77 ( .A(aes_core_sbox_inst_n196), .Y(
        aes_core_sbox_inst_n201) );
  INVX1 aes_core_sbox_inst_U76 ( .A(aes_core_sbox_inst_n156), .Y(
        aes_core_sbox_inst_n162) );
  OR2X2 aes_core_sbox_inst_U75 ( .A(aes_core_sbox_inst_n46), .B(
        aes_core_sbox_inst_n43), .Y(aes_core_sbox_inst_n2) );
  INVX1 aes_core_sbox_inst_U74 ( .A(aes_core_n7), .Y(aes_core_sbox_inst_n190)
         );
  INVX1 aes_core_sbox_inst_U73 ( .A(aes_core_n27), .Y(aes_core_sbox_inst_n153)
         );
  NOR2X1 aes_core_sbox_inst_U72 ( .A(aes_core_sbox_inst_n201), .B(
        aes_core_sbox_inst_n195), .Y(aes_core_sbox_inst_n384) );
  INVX1 aes_core_sbox_inst_U71 ( .A(aes_core_n27), .Y(aes_core_sbox_inst_n155)
         );
  INVX1 aes_core_sbox_inst_U70 ( .A(aes_core_n31), .Y(aes_core_sbox_inst_n149)
         );
  INVX1 aes_core_sbox_inst_U69 ( .A(aes_core_n3), .Y(aes_core_sbox_inst_n195)
         );
  OR2X2 aes_core_sbox_inst_U68 ( .A(aes_core_sbox_inst_n162), .B(
        aes_core_sbox_inst_n153), .Y(aes_core_sbox_inst_n1) );
  CLKINVX3 aes_core_sbox_inst_U67 ( .A(aes_core_sbox_inst_n178), .Y(
        aes_core_sbox_inst_n174) );
  INVX1 aes_core_sbox_inst_U66 ( .A(aes_core_n19), .Y(aes_core_sbox_inst_n173)
         );
  INVX1 aes_core_sbox_inst_U65 ( .A(aes_core_n23), .Y(aes_core_sbox_inst_n168)
         );
  INVX2 aes_core_sbox_inst_U64 ( .A(aes_core_sbox_inst_n150), .Y(
        aes_core_sbox_inst_n146) );
  INVX1 aes_core_sbox_inst_U63 ( .A(aes_core_sbox_inst_n551), .Y(
        aes_core_sbox_inst_n1688) );
  NOR4BX1 aes_core_sbox_inst_U62 ( .AN(aes_core_sbox_inst_n645), .B(
        aes_core_sbox_inst_n646), .C(aes_core_sbox_inst_n647), .D(
        aes_core_sbox_inst_n648), .Y(aes_core_sbox_inst_n605) );
  AOI211X1 aes_core_sbox_inst_U61 ( .A0(aes_core_sbox_inst_n607), .A1(
        aes_core_sbox_inst_n608), .B0(aes_core_sbox_inst_n609), .C0(
        aes_core_sbox_inst_n610), .Y(aes_core_sbox_inst_n606) );
  NOR3BX1 aes_core_sbox_inst_U60 ( .AN(aes_core_sbox_inst_n659), .B(
        aes_core_sbox_inst_n660), .C(aes_core_sbox_inst_n661), .Y(
        aes_core_sbox_inst_n604) );
  OAI222X4 aes_core_sbox_inst_U59 ( .A0(aes_core_sbox_inst_n604), .A1(
        aes_core_sbox_inst_n204), .B0(aes_core_sbox_inst_n605), .B1(
        aes_core_sbox_inst_n205), .C0(aes_core_n33), .C1(
        aes_core_sbox_inst_n606), .Y(aes_core_new_sboxw[31]) );
  NOR2X2 aes_core_sbox_inst_U58 ( .A(aes_core_sbox_inst_n55), .B(
        aes_core_sbox_inst_n186), .Y(aes_core_sbox_inst_n404) );
  NOR2X2 aes_core_sbox_inst_U57 ( .A(aes_core_sbox_inst_n60), .B(
        aes_core_sbox_inst_n164), .Y(aes_core_sbox_inst_n999) );
  AOI222X1 aes_core_sbox_inst_U56 ( .A0(aes_core_sbox_inst_n64), .A1(
        aes_core_sbox_inst_n795), .B0(aes_core_sbox_inst_n796), .B1(
        aes_core_sbox_inst_n797), .C0(aes_core_sbox_inst_n673), .C1(
        aes_core_sbox_inst_n798), .Y(aes_core_sbox_inst_n794) );
  AOI211X1 aes_core_sbox_inst_U55 ( .A0(aes_core_sbox_inst_n64), .A1(
        aes_core_sbox_inst_n814), .B0(aes_core_sbox_inst_n212), .C0(
        aes_core_sbox_inst_n815), .Y(aes_core_sbox_inst_n793) );
  OAI22X2 aes_core_sbox_inst_U54 ( .A0(aes_core_n33), .A1(
        aes_core_sbox_inst_n793), .B0(aes_core_sbox_inst_n794), .B1(
        aes_core_sbox_inst_n206), .Y(aes_core_new_sboxw[28]) );
  AOI211X1 aes_core_sbox_inst_U53 ( .A0(aes_core_sbox_inst_n832), .A1(
        aes_core_sbox_inst_n833), .B0(aes_core_sbox_inst_n834), .C0(
        aes_core_sbox_inst_n835), .Y(aes_core_sbox_inst_n831) );
  CLKINVX3 aes_core_sbox_inst_U52 ( .A(aes_core_sbox_inst_n831), .Y(
        aes_core_new_sboxw[27]) );
  BUFX12 aes_core_sbox_inst_U51 ( .A(aes_core_sbox_inst_n1672), .Y(
        aes_core_sbox_inst_n38) );
  NOR2X2 aes_core_sbox_inst_U50 ( .A(aes_core_sbox_inst_n42), .B(
        aes_core_sbox_inst_n57), .Y(aes_core_sbox_inst_n281) );
  BUFX8 aes_core_sbox_inst_U49 ( .A(aes_core_sbox_inst_n281), .Y(
        aes_core_sbox_inst_n79) );
  NOR2X2 aes_core_sbox_inst_U48 ( .A(aes_core_sbox_inst_n1651), .B(
        aes_core_sbox_inst_n43), .Y(aes_core_sbox_inst_n1355) );
  BUFX4 aes_core_sbox_inst_U47 ( .A(aes_core_n10), .Y(aes_core_sbox_inst_n57)
         );
  BUFX4 aes_core_sbox_inst_U46 ( .A(aes_core_n12), .Y(aes_core_sbox_inst_n59)
         );
  BUFX8 aes_core_sbox_inst_U45 ( .A(aes_core_sbox_inst_n1029), .Y(
        aes_core_sbox_inst_n104) );
  CLKBUFX8 aes_core_sbox_inst_U44 ( .A(aes_core_sbox_inst_n1595), .Y(
        aes_core_sbox_inst_n23) );
  NOR2X2 aes_core_sbox_inst_U43 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_sbox_inst_n1594), .Y(aes_core_sbox_inst_n1004) );
  CLKBUFX8 aes_core_sbox_inst_U42 ( .A(aes_core_sbox_inst_n1004), .Y(
        aes_core_sbox_inst_n94) );
  BUFX12 aes_core_sbox_inst_U41 ( .A(aes_core_sbox_inst_n981), .Y(
        aes_core_sbox_inst_n96) );
  NOR2X1 aes_core_sbox_inst_U40 ( .A(aes_core_sbox_inst_n26), .B(
        aes_core_sbox_inst_n165), .Y(aes_core_sbox_inst_n994) );
  NOR2X1 aes_core_sbox_inst_U39 ( .A(aes_core_sbox_inst_n590), .B(aes_core_n6), 
        .Y(aes_core_sbox_inst_n446) );
  CLKBUFX8 aes_core_sbox_inst_U38 ( .A(aes_core_sbox_inst_n1713), .Y(
        aes_core_sbox_inst_n49) );
  NOR2X2 aes_core_sbox_inst_U37 ( .A(aes_core_sbox_inst_n138), .B(
        aes_core_sbox_inst_n69), .Y(aes_core_sbox_inst_n386) );
  CLKBUFX8 aes_core_sbox_inst_U36 ( .A(aes_core_sbox_inst_n386), .Y(
        aes_core_sbox_inst_n70) );
  BUFX4 aes_core_sbox_inst_U35 ( .A(aes_core_sbox_inst_n1670), .Y(
        aes_core_sbox_inst_n37) );
  BUFX3 aes_core_sbox_inst_U34 ( .A(aes_core_sbox_inst_n274), .Y(
        aes_core_sbox_inst_n88) );
  INVX1 aes_core_sbox_inst_U33 ( .A(aes_core_sbox_inst_n112), .Y(
        aes_core_sbox_inst_n229) );
  CLKINVX3 aes_core_sbox_inst_U32 ( .A(aes_core_sbox_inst_n77), .Y(
        aes_core_sbox_inst_n1724) );
  CLKINVX3 aes_core_sbox_inst_U31 ( .A(aes_core_sbox_inst_n83), .Y(
        aes_core_sbox_inst_n1661) );
  INVX4 aes_core_sbox_inst_U30 ( .A(aes_core_sbox_inst_n82), .Y(
        aes_core_sbox_inst_n1663) );
  INVX4 aes_core_sbox_inst_U29 ( .A(aes_core_sbox_inst_n66), .Y(
        aes_core_sbox_inst_n1703) );
  CLKINVX3 aes_core_sbox_inst_U28 ( .A(aes_core_sbox_inst_n103), .Y(
        aes_core_sbox_inst_n1606) );
  INVX4 aes_core_sbox_inst_U27 ( .A(aes_core_sbox_inst_n101), .Y(
        aes_core_sbox_inst_n1584) );
  CLKBUFX8 aes_core_sbox_inst_U26 ( .A(aes_core_sbox_inst_n1585), .Y(
        aes_core_sbox_inst_n22) );
  NOR2X1 aes_core_sbox_inst_U25 ( .A(aes_core_sbox_inst_n1579), .B(
        aes_core_sbox_inst_n25), .Y(aes_core_sbox_inst_n1198) );
  INVX1 aes_core_sbox_inst_U24 ( .A(aes_core_sbox_inst_n3), .Y(
        aes_core_sbox_inst_n1700) );
  INVX2 aes_core_sbox_inst_U23 ( .A(aes_core_sbox_inst_n1045), .Y(
        aes_core_sbox_inst_n1582) );
  CLKINVX3 aes_core_sbox_inst_U22 ( .A(aes_core_sbox_inst_n91), .Y(
        aes_core_sbox_inst_n1594) );
  NOR2X1 aes_core_sbox_inst_U21 ( .A(aes_core_sbox_inst_n191), .B(
        aes_core_sbox_inst_n199), .Y(aes_core_sbox_inst_n437) );
  NOR2X2 aes_core_sbox_inst_U20 ( .A(aes_core_sbox_inst_n857), .B(aes_core_n30), .Y(aes_core_sbox_inst_n679) );
  CLKBUFX8 aes_core_sbox_inst_U19 ( .A(aes_core_sbox_inst_n635), .Y(
        aes_core_sbox_inst_n105) );
  NOR2X1 aes_core_sbox_inst_U18 ( .A(aes_core_sbox_inst_n16), .B(
        aes_core_sbox_inst_n19), .Y(aes_core_sbox_inst_n710) );
  CLKINVX3 aes_core_sbox_inst_U17 ( .A(aes_core_sbox_inst_n110), .Y(
        aes_core_sbox_inst_n243) );
  NOR2X1 aes_core_sbox_inst_U16 ( .A(aes_core_sbox_inst_n163), .B(
        aes_core_sbox_inst_n151), .Y(aes_core_sbox_inst_n9) );
  CLKBUFX8 aes_core_sbox_inst_U15 ( .A(aes_core_sbox_inst_n642), .Y(
        aes_core_sbox_inst_n108) );
  CLKINVX3 aes_core_sbox_inst_U14 ( .A(aes_core_sbox_inst_n632), .Y(
        aes_core_sbox_inst_n221) );
  NOR2X1 aes_core_sbox_inst_U13 ( .A(aes_core_sbox_inst_n145), .B(
        aes_core_sbox_inst_n1654), .Y(aes_core_sbox_inst_n1498) );
  CLKINVX3 aes_core_sbox_inst_U12 ( .A(aes_core_sbox_inst_n115), .Y(
        aes_core_sbox_inst_n247) );
  NOR2X2 aes_core_sbox_inst_U11 ( .A(aes_core_sbox_inst_n51), .B(aes_core_n5), 
        .Y(aes_core_sbox_inst_n561) );
  INVX1 aes_core_sbox_inst_U10 ( .A(aes_core_sbox_inst_n469), .Y(
        aes_core_sbox_inst_n1698) );
  INVX1 aes_core_sbox_inst_U9 ( .A(aes_core_sbox_inst_n106), .Y(
        aes_core_sbox_inst_n226) );
  BUFX3 aes_core_sbox_inst_U8 ( .A(aes_core_sbox_inst_n226), .Y(
        aes_core_sbox_inst_n14) );
  INVX1 aes_core_sbox_inst_U7 ( .A(aes_core_sbox_inst_n703), .Y(
        aes_core_sbox_inst_n230) );
  NOR2X1 aes_core_sbox_inst_U6 ( .A(aes_core_sbox_inst_n117), .B(
        aes_core_sbox_inst_n16), .Y(aes_core_sbox_inst_n791) );
  INVX1 aes_core_sbox_inst_U5 ( .A(aes_core_sbox_inst_n947), .Y(
        aes_core_sbox_inst_n219) );
  NOR2X1 aes_core_sbox_inst_U4 ( .A(aes_core_sbox_inst_n34), .B(
        aes_core_sbox_inst_n38), .Y(aes_core_sbox_inst_n305) );
  INVX4 aes_core_sbox_inst_U3 ( .A(aes_core_sbox_inst_n72), .Y(
        aes_core_sbox_inst_n1718) );
  AOI21X1 aes_core_sbox_inst_U2 ( .A0(aes_core_sbox_inst_n115), .A1(
        aes_core_sbox_inst_n152), .B0(aes_core_sbox_inst_n718), .Y(
        aes_core_sbox_inst_n716) );
  OAI22X1 aes_core_sbox_inst_U1 ( .A0(aes_core_sbox_inst_n146), .A1(
        aes_core_sbox_inst_n715), .B0(aes_core_sbox_inst_n716), .B1(
        aes_core_sbox_inst_n148), .Y(aes_core_sbox_inst_n714) );
  INVX1 reg_in_U1034 ( .A(reg_in_plain_text[255]), .Y(reg_in_n808) );
  INVX1 reg_in_U1033 ( .A(reg_in_plain_text[254]), .Y(reg_in_n840) );
  INVX1 reg_in_U1032 ( .A(reg_in_plain_text[253]), .Y(reg_in_n872) );
  INVX1 reg_in_U1031 ( .A(reg_in_plain_text[252]), .Y(reg_in_n904) );
  INVX1 reg_in_U1030 ( .A(reg_in_plain_text[251]), .Y(reg_in_n936) );
  INVX1 reg_in_U1029 ( .A(reg_in_plain_text[250]), .Y(reg_in_n968) );
  INVX1 reg_in_U1028 ( .A(reg_in_plain_text[249]), .Y(reg_in_n1000) );
  INVX1 reg_in_U1027 ( .A(reg_in_plain_text[248]), .Y(reg_in_n1032) );
  INVX1 reg_in_U1026 ( .A(reg_in_plain_text[15]), .Y(reg_in_n778) );
  INVX1 reg_in_U1025 ( .A(reg_in_plain_text[23]), .Y(reg_in_n779) );
  INVX1 reg_in_U1024 ( .A(reg_in_plain_text[31]), .Y(reg_in_n780) );
  INVX1 reg_in_U1023 ( .A(reg_in_plain_text[39]), .Y(reg_in_n781) );
  INVX1 reg_in_U1022 ( .A(reg_in_plain_text[47]), .Y(reg_in_n782) );
  INVX1 reg_in_U1021 ( .A(reg_in_plain_text[55]), .Y(reg_in_n783) );
  INVX1 reg_in_U1020 ( .A(reg_in_plain_text[63]), .Y(reg_in_n784) );
  INVX1 reg_in_U1019 ( .A(reg_in_plain_text[71]), .Y(reg_in_n785) );
  INVX1 reg_in_U1018 ( .A(reg_in_plain_text[79]), .Y(reg_in_n786) );
  INVX1 reg_in_U1017 ( .A(reg_in_plain_text[87]), .Y(reg_in_n787) );
  INVX1 reg_in_U1016 ( .A(reg_in_plain_text[95]), .Y(reg_in_n788) );
  INVX1 reg_in_U1015 ( .A(reg_in_plain_text[103]), .Y(reg_in_n789) );
  INVX1 reg_in_U1014 ( .A(reg_in_plain_text[111]), .Y(reg_in_n790) );
  INVX1 reg_in_U1013 ( .A(reg_in_plain_text[119]), .Y(reg_in_n791) );
  INVX1 reg_in_U1012 ( .A(reg_in_plain_text[127]), .Y(reg_in_n792) );
  INVX1 reg_in_U1011 ( .A(reg_in_plain_text[135]), .Y(reg_in_n793) );
  INVX1 reg_in_U1010 ( .A(reg_in_plain_text[143]), .Y(reg_in_n794) );
  INVX1 reg_in_U1009 ( .A(reg_in_plain_text[151]), .Y(reg_in_n795) );
  INVX1 reg_in_U1008 ( .A(reg_in_plain_text[159]), .Y(reg_in_n796) );
  INVX1 reg_in_U1007 ( .A(reg_in_plain_text[167]), .Y(reg_in_n797) );
  INVX1 reg_in_U1006 ( .A(reg_in_plain_text[175]), .Y(reg_in_n798) );
  INVX1 reg_in_U1005 ( .A(reg_in_plain_text[183]), .Y(reg_in_n799) );
  INVX1 reg_in_U1004 ( .A(reg_in_plain_text[191]), .Y(reg_in_n800) );
  INVX1 reg_in_U1003 ( .A(reg_in_plain_text[199]), .Y(reg_in_n801) );
  INVX1 reg_in_U1002 ( .A(reg_in_plain_text[207]), .Y(reg_in_n802) );
  INVX1 reg_in_U1001 ( .A(reg_in_plain_text[215]), .Y(reg_in_n803) );
  INVX1 reg_in_U1000 ( .A(reg_in_plain_text[223]), .Y(reg_in_n804) );
  INVX1 reg_in_U999 ( .A(reg_in_plain_text[231]), .Y(reg_in_n805) );
  INVX1 reg_in_U998 ( .A(reg_in_plain_text[239]), .Y(reg_in_n806) );
  INVX1 reg_in_U997 ( .A(reg_in_plain_text[247]), .Y(reg_in_n807) );
  INVX1 reg_in_U996 ( .A(reg_in_plain_text[14]), .Y(reg_in_n810) );
  INVX1 reg_in_U995 ( .A(reg_in_plain_text[22]), .Y(reg_in_n811) );
  INVX1 reg_in_U994 ( .A(reg_in_plain_text[30]), .Y(reg_in_n812) );
  INVX1 reg_in_U993 ( .A(reg_in_plain_text[38]), .Y(reg_in_n813) );
  INVX1 reg_in_U992 ( .A(reg_in_plain_text[46]), .Y(reg_in_n814) );
  INVX1 reg_in_U991 ( .A(reg_in_plain_text[54]), .Y(reg_in_n815) );
  INVX1 reg_in_U990 ( .A(reg_in_plain_text[62]), .Y(reg_in_n816) );
  INVX1 reg_in_U989 ( .A(reg_in_plain_text[70]), .Y(reg_in_n817) );
  INVX1 reg_in_U988 ( .A(reg_in_plain_text[78]), .Y(reg_in_n818) );
  INVX1 reg_in_U987 ( .A(reg_in_plain_text[86]), .Y(reg_in_n819) );
  INVX1 reg_in_U986 ( .A(reg_in_plain_text[94]), .Y(reg_in_n820) );
  INVX1 reg_in_U985 ( .A(reg_in_plain_text[102]), .Y(reg_in_n821) );
  INVX1 reg_in_U984 ( .A(reg_in_plain_text[110]), .Y(reg_in_n822) );
  INVX1 reg_in_U983 ( .A(reg_in_plain_text[118]), .Y(reg_in_n823) );
  INVX1 reg_in_U982 ( .A(reg_in_plain_text[126]), .Y(reg_in_n824) );
  INVX1 reg_in_U981 ( .A(reg_in_plain_text[134]), .Y(reg_in_n825) );
  INVX1 reg_in_U980 ( .A(reg_in_plain_text[142]), .Y(reg_in_n826) );
  INVX1 reg_in_U979 ( .A(reg_in_plain_text[150]), .Y(reg_in_n827) );
  INVX1 reg_in_U978 ( .A(reg_in_plain_text[158]), .Y(reg_in_n828) );
  INVX1 reg_in_U977 ( .A(reg_in_plain_text[166]), .Y(reg_in_n829) );
  INVX1 reg_in_U976 ( .A(reg_in_plain_text[174]), .Y(reg_in_n830) );
  INVX1 reg_in_U975 ( .A(reg_in_plain_text[182]), .Y(reg_in_n831) );
  INVX1 reg_in_U974 ( .A(reg_in_plain_text[190]), .Y(reg_in_n832) );
  INVX1 reg_in_U973 ( .A(reg_in_plain_text[198]), .Y(reg_in_n833) );
  INVX1 reg_in_U972 ( .A(reg_in_plain_text[206]), .Y(reg_in_n834) );
  INVX1 reg_in_U971 ( .A(reg_in_plain_text[214]), .Y(reg_in_n835) );
  INVX1 reg_in_U970 ( .A(reg_in_plain_text[222]), .Y(reg_in_n836) );
  INVX1 reg_in_U969 ( .A(reg_in_plain_text[230]), .Y(reg_in_n837) );
  INVX1 reg_in_U968 ( .A(reg_in_plain_text[238]), .Y(reg_in_n838) );
  INVX1 reg_in_U967 ( .A(reg_in_plain_text[246]), .Y(reg_in_n839) );
  INVX1 reg_in_U966 ( .A(reg_in_plain_text[13]), .Y(reg_in_n842) );
  INVX1 reg_in_U965 ( .A(reg_in_plain_text[21]), .Y(reg_in_n843) );
  INVX1 reg_in_U964 ( .A(reg_in_plain_text[29]), .Y(reg_in_n844) );
  INVX1 reg_in_U963 ( .A(reg_in_plain_text[37]), .Y(reg_in_n845) );
  INVX1 reg_in_U962 ( .A(reg_in_plain_text[45]), .Y(reg_in_n846) );
  INVX1 reg_in_U961 ( .A(reg_in_plain_text[53]), .Y(reg_in_n847) );
  INVX1 reg_in_U960 ( .A(reg_in_plain_text[61]), .Y(reg_in_n848) );
  INVX1 reg_in_U959 ( .A(reg_in_plain_text[69]), .Y(reg_in_n849) );
  INVX1 reg_in_U958 ( .A(reg_in_plain_text[77]), .Y(reg_in_n850) );
  INVX1 reg_in_U957 ( .A(reg_in_plain_text[85]), .Y(reg_in_n851) );
  INVX1 reg_in_U956 ( .A(reg_in_plain_text[93]), .Y(reg_in_n852) );
  INVX1 reg_in_U955 ( .A(reg_in_plain_text[101]), .Y(reg_in_n853) );
  INVX1 reg_in_U954 ( .A(reg_in_plain_text[109]), .Y(reg_in_n854) );
  INVX1 reg_in_U953 ( .A(reg_in_plain_text[117]), .Y(reg_in_n855) );
  INVX1 reg_in_U952 ( .A(reg_in_plain_text[125]), .Y(reg_in_n856) );
  INVX1 reg_in_U951 ( .A(reg_in_plain_text[133]), .Y(reg_in_n857) );
  INVX1 reg_in_U950 ( .A(reg_in_plain_text[141]), .Y(reg_in_n858) );
  INVX1 reg_in_U949 ( .A(reg_in_plain_text[149]), .Y(reg_in_n859) );
  INVX1 reg_in_U948 ( .A(reg_in_plain_text[157]), .Y(reg_in_n860) );
  INVX1 reg_in_U947 ( .A(reg_in_plain_text[165]), .Y(reg_in_n861) );
  INVX1 reg_in_U946 ( .A(reg_in_plain_text[173]), .Y(reg_in_n862) );
  INVX1 reg_in_U945 ( .A(reg_in_plain_text[181]), .Y(reg_in_n863) );
  INVX1 reg_in_U944 ( .A(reg_in_plain_text[189]), .Y(reg_in_n864) );
  INVX1 reg_in_U943 ( .A(reg_in_plain_text[197]), .Y(reg_in_n865) );
  INVX1 reg_in_U942 ( .A(reg_in_plain_text[205]), .Y(reg_in_n866) );
  INVX1 reg_in_U941 ( .A(reg_in_plain_text[213]), .Y(reg_in_n867) );
  INVX1 reg_in_U940 ( .A(reg_in_plain_text[221]), .Y(reg_in_n868) );
  INVX1 reg_in_U939 ( .A(reg_in_plain_text[229]), .Y(reg_in_n869) );
  INVX1 reg_in_U938 ( .A(reg_in_plain_text[237]), .Y(reg_in_n870) );
  INVX1 reg_in_U937 ( .A(reg_in_plain_text[245]), .Y(reg_in_n871) );
  INVX1 reg_in_U936 ( .A(reg_in_plain_text[12]), .Y(reg_in_n874) );
  INVX1 reg_in_U935 ( .A(reg_in_plain_text[20]), .Y(reg_in_n875) );
  INVX1 reg_in_U934 ( .A(reg_in_plain_text[28]), .Y(reg_in_n876) );
  INVX1 reg_in_U933 ( .A(reg_in_plain_text[36]), .Y(reg_in_n877) );
  INVX1 reg_in_U932 ( .A(reg_in_plain_text[44]), .Y(reg_in_n878) );
  INVX1 reg_in_U931 ( .A(reg_in_plain_text[52]), .Y(reg_in_n879) );
  INVX1 reg_in_U930 ( .A(reg_in_plain_text[60]), .Y(reg_in_n880) );
  INVX1 reg_in_U929 ( .A(reg_in_plain_text[68]), .Y(reg_in_n881) );
  INVX1 reg_in_U928 ( .A(reg_in_plain_text[76]), .Y(reg_in_n882) );
  INVX1 reg_in_U927 ( .A(reg_in_plain_text[84]), .Y(reg_in_n883) );
  INVX1 reg_in_U926 ( .A(reg_in_plain_text[92]), .Y(reg_in_n884) );
  INVX1 reg_in_U925 ( .A(reg_in_plain_text[100]), .Y(reg_in_n885) );
  INVX1 reg_in_U924 ( .A(reg_in_plain_text[108]), .Y(reg_in_n886) );
  INVX1 reg_in_U923 ( .A(reg_in_plain_text[116]), .Y(reg_in_n887) );
  INVX1 reg_in_U922 ( .A(reg_in_plain_text[124]), .Y(reg_in_n888) );
  INVX1 reg_in_U921 ( .A(reg_in_plain_text[132]), .Y(reg_in_n889) );
  INVX1 reg_in_U920 ( .A(reg_in_plain_text[140]), .Y(reg_in_n890) );
  INVX1 reg_in_U919 ( .A(reg_in_plain_text[148]), .Y(reg_in_n891) );
  INVX1 reg_in_U918 ( .A(reg_in_plain_text[156]), .Y(reg_in_n892) );
  INVX1 reg_in_U917 ( .A(reg_in_plain_text[164]), .Y(reg_in_n893) );
  INVX1 reg_in_U916 ( .A(reg_in_plain_text[172]), .Y(reg_in_n894) );
  INVX1 reg_in_U915 ( .A(reg_in_plain_text[180]), .Y(reg_in_n895) );
  INVX1 reg_in_U914 ( .A(reg_in_plain_text[188]), .Y(reg_in_n896) );
  INVX1 reg_in_U913 ( .A(reg_in_plain_text[196]), .Y(reg_in_n897) );
  INVX1 reg_in_U912 ( .A(reg_in_plain_text[204]), .Y(reg_in_n898) );
  INVX1 reg_in_U911 ( .A(reg_in_plain_text[212]), .Y(reg_in_n899) );
  INVX1 reg_in_U910 ( .A(reg_in_plain_text[220]), .Y(reg_in_n900) );
  INVX1 reg_in_U909 ( .A(reg_in_plain_text[228]), .Y(reg_in_n901) );
  INVX1 reg_in_U908 ( .A(reg_in_plain_text[236]), .Y(reg_in_n902) );
  INVX1 reg_in_U907 ( .A(reg_in_plain_text[244]), .Y(reg_in_n903) );
  INVX1 reg_in_U906 ( .A(reg_in_plain_text[11]), .Y(reg_in_n906) );
  INVX1 reg_in_U905 ( .A(reg_in_plain_text[19]), .Y(reg_in_n907) );
  INVX1 reg_in_U904 ( .A(reg_in_plain_text[27]), .Y(reg_in_n908) );
  INVX1 reg_in_U903 ( .A(reg_in_plain_text[35]), .Y(reg_in_n909) );
  INVX1 reg_in_U902 ( .A(reg_in_plain_text[43]), .Y(reg_in_n910) );
  INVX1 reg_in_U901 ( .A(reg_in_plain_text[51]), .Y(reg_in_n911) );
  INVX1 reg_in_U900 ( .A(reg_in_plain_text[59]), .Y(reg_in_n912) );
  INVX1 reg_in_U899 ( .A(reg_in_plain_text[67]), .Y(reg_in_n913) );
  INVX1 reg_in_U898 ( .A(reg_in_plain_text[75]), .Y(reg_in_n914) );
  INVX1 reg_in_U897 ( .A(reg_in_plain_text[83]), .Y(reg_in_n915) );
  INVX1 reg_in_U896 ( .A(reg_in_plain_text[91]), .Y(reg_in_n916) );
  INVX1 reg_in_U895 ( .A(reg_in_plain_text[99]), .Y(reg_in_n917) );
  INVX1 reg_in_U894 ( .A(reg_in_plain_text[107]), .Y(reg_in_n918) );
  INVX1 reg_in_U893 ( .A(reg_in_plain_text[115]), .Y(reg_in_n919) );
  INVX1 reg_in_U892 ( .A(reg_in_plain_text[123]), .Y(reg_in_n920) );
  INVX1 reg_in_U891 ( .A(reg_in_plain_text[131]), .Y(reg_in_n921) );
  INVX1 reg_in_U890 ( .A(reg_in_plain_text[139]), .Y(reg_in_n922) );
  INVX1 reg_in_U889 ( .A(reg_in_plain_text[147]), .Y(reg_in_n923) );
  INVX1 reg_in_U888 ( .A(reg_in_plain_text[155]), .Y(reg_in_n924) );
  INVX1 reg_in_U887 ( .A(reg_in_plain_text[163]), .Y(reg_in_n925) );
  INVX1 reg_in_U886 ( .A(reg_in_plain_text[171]), .Y(reg_in_n926) );
  INVX1 reg_in_U885 ( .A(reg_in_plain_text[179]), .Y(reg_in_n927) );
  INVX1 reg_in_U884 ( .A(reg_in_plain_text[187]), .Y(reg_in_n928) );
  INVX1 reg_in_U883 ( .A(reg_in_plain_text[195]), .Y(reg_in_n929) );
  INVX1 reg_in_U882 ( .A(reg_in_plain_text[203]), .Y(reg_in_n930) );
  INVX1 reg_in_U881 ( .A(reg_in_plain_text[211]), .Y(reg_in_n931) );
  INVX1 reg_in_U880 ( .A(reg_in_plain_text[219]), .Y(reg_in_n932) );
  INVX1 reg_in_U879 ( .A(reg_in_plain_text[227]), .Y(reg_in_n933) );
  INVX1 reg_in_U878 ( .A(reg_in_plain_text[235]), .Y(reg_in_n934) );
  INVX1 reg_in_U877 ( .A(reg_in_plain_text[243]), .Y(reg_in_n935) );
  INVX1 reg_in_U876 ( .A(reg_in_plain_text[10]), .Y(reg_in_n938) );
  INVX1 reg_in_U875 ( .A(reg_in_plain_text[18]), .Y(reg_in_n939) );
  INVX1 reg_in_U874 ( .A(reg_in_plain_text[26]), .Y(reg_in_n940) );
  INVX1 reg_in_U873 ( .A(reg_in_plain_text[34]), .Y(reg_in_n941) );
  INVX1 reg_in_U872 ( .A(reg_in_plain_text[42]), .Y(reg_in_n942) );
  INVX1 reg_in_U871 ( .A(reg_in_plain_text[50]), .Y(reg_in_n943) );
  INVX1 reg_in_U870 ( .A(reg_in_plain_text[58]), .Y(reg_in_n944) );
  INVX1 reg_in_U869 ( .A(reg_in_plain_text[66]), .Y(reg_in_n945) );
  INVX1 reg_in_U868 ( .A(reg_in_plain_text[74]), .Y(reg_in_n946) );
  INVX1 reg_in_U867 ( .A(reg_in_plain_text[82]), .Y(reg_in_n947) );
  INVX1 reg_in_U866 ( .A(reg_in_plain_text[90]), .Y(reg_in_n948) );
  INVX1 reg_in_U865 ( .A(reg_in_plain_text[98]), .Y(reg_in_n949) );
  INVX1 reg_in_U864 ( .A(reg_in_plain_text[106]), .Y(reg_in_n950) );
  INVX1 reg_in_U863 ( .A(reg_in_plain_text[114]), .Y(reg_in_n951) );
  INVX1 reg_in_U862 ( .A(reg_in_plain_text[122]), .Y(reg_in_n952) );
  INVX1 reg_in_U861 ( .A(reg_in_plain_text[130]), .Y(reg_in_n953) );
  INVX1 reg_in_U860 ( .A(reg_in_plain_text[138]), .Y(reg_in_n954) );
  INVX1 reg_in_U859 ( .A(reg_in_plain_text[146]), .Y(reg_in_n955) );
  INVX1 reg_in_U858 ( .A(reg_in_plain_text[154]), .Y(reg_in_n956) );
  INVX1 reg_in_U857 ( .A(reg_in_plain_text[162]), .Y(reg_in_n957) );
  INVX1 reg_in_U856 ( .A(reg_in_plain_text[170]), .Y(reg_in_n958) );
  INVX1 reg_in_U855 ( .A(reg_in_plain_text[178]), .Y(reg_in_n959) );
  INVX1 reg_in_U854 ( .A(reg_in_plain_text[186]), .Y(reg_in_n960) );
  INVX1 reg_in_U853 ( .A(reg_in_plain_text[194]), .Y(reg_in_n961) );
  INVX1 reg_in_U852 ( .A(reg_in_plain_text[202]), .Y(reg_in_n962) );
  INVX1 reg_in_U851 ( .A(reg_in_plain_text[210]), .Y(reg_in_n963) );
  INVX1 reg_in_U850 ( .A(reg_in_plain_text[218]), .Y(reg_in_n964) );
  INVX1 reg_in_U849 ( .A(reg_in_plain_text[226]), .Y(reg_in_n965) );
  INVX1 reg_in_U848 ( .A(reg_in_plain_text[234]), .Y(reg_in_n966) );
  INVX1 reg_in_U847 ( .A(reg_in_plain_text[242]), .Y(reg_in_n967) );
  INVX1 reg_in_U846 ( .A(reg_in_plain_text[9]), .Y(reg_in_n970) );
  INVX1 reg_in_U845 ( .A(reg_in_plain_text[17]), .Y(reg_in_n971) );
  INVX1 reg_in_U844 ( .A(reg_in_plain_text[25]), .Y(reg_in_n972) );
  INVX1 reg_in_U843 ( .A(reg_in_plain_text[33]), .Y(reg_in_n973) );
  INVX1 reg_in_U842 ( .A(reg_in_plain_text[41]), .Y(reg_in_n974) );
  INVX1 reg_in_U841 ( .A(reg_in_plain_text[49]), .Y(reg_in_n975) );
  INVX1 reg_in_U840 ( .A(reg_in_plain_text[57]), .Y(reg_in_n976) );
  INVX1 reg_in_U839 ( .A(reg_in_plain_text[65]), .Y(reg_in_n977) );
  INVX1 reg_in_U838 ( .A(reg_in_plain_text[73]), .Y(reg_in_n978) );
  INVX1 reg_in_U837 ( .A(reg_in_plain_text[81]), .Y(reg_in_n979) );
  INVX1 reg_in_U836 ( .A(reg_in_plain_text[89]), .Y(reg_in_n980) );
  INVX1 reg_in_U835 ( .A(reg_in_plain_text[97]), .Y(reg_in_n981) );
  INVX1 reg_in_U834 ( .A(reg_in_plain_text[105]), .Y(reg_in_n982) );
  INVX1 reg_in_U833 ( .A(reg_in_plain_text[113]), .Y(reg_in_n983) );
  INVX1 reg_in_U832 ( .A(reg_in_plain_text[121]), .Y(reg_in_n984) );
  INVX1 reg_in_U831 ( .A(reg_in_plain_text[129]), .Y(reg_in_n985) );
  INVX1 reg_in_U830 ( .A(reg_in_plain_text[137]), .Y(reg_in_n986) );
  INVX1 reg_in_U829 ( .A(reg_in_plain_text[145]), .Y(reg_in_n987) );
  INVX1 reg_in_U828 ( .A(reg_in_plain_text[153]), .Y(reg_in_n988) );
  INVX1 reg_in_U827 ( .A(reg_in_plain_text[161]), .Y(reg_in_n989) );
  INVX1 reg_in_U826 ( .A(reg_in_plain_text[169]), .Y(reg_in_n990) );
  INVX1 reg_in_U825 ( .A(reg_in_plain_text[177]), .Y(reg_in_n991) );
  INVX1 reg_in_U824 ( .A(reg_in_plain_text[185]), .Y(reg_in_n992) );
  INVX1 reg_in_U823 ( .A(reg_in_plain_text[193]), .Y(reg_in_n993) );
  INVX1 reg_in_U822 ( .A(reg_in_plain_text[201]), .Y(reg_in_n994) );
  INVX1 reg_in_U821 ( .A(reg_in_plain_text[209]), .Y(reg_in_n995) );
  INVX1 reg_in_U820 ( .A(reg_in_plain_text[217]), .Y(reg_in_n996) );
  INVX1 reg_in_U819 ( .A(reg_in_plain_text[225]), .Y(reg_in_n997) );
  INVX1 reg_in_U818 ( .A(reg_in_plain_text[233]), .Y(reg_in_n998) );
  INVX1 reg_in_U817 ( .A(reg_in_plain_text[241]), .Y(reg_in_n999) );
  INVX1 reg_in_U816 ( .A(reg_in_plain_text[8]), .Y(reg_in_n1002) );
  INVX1 reg_in_U815 ( .A(reg_in_plain_text[16]), .Y(reg_in_n1003) );
  INVX1 reg_in_U814 ( .A(reg_in_plain_text[24]), .Y(reg_in_n1004) );
  INVX1 reg_in_U813 ( .A(reg_in_plain_text[32]), .Y(reg_in_n1005) );
  INVX1 reg_in_U812 ( .A(reg_in_plain_text[40]), .Y(reg_in_n1006) );
  INVX1 reg_in_U811 ( .A(reg_in_plain_text[48]), .Y(reg_in_n1007) );
  INVX1 reg_in_U810 ( .A(reg_in_plain_text[56]), .Y(reg_in_n1008) );
  INVX1 reg_in_U809 ( .A(reg_in_plain_text[64]), .Y(reg_in_n1009) );
  INVX1 reg_in_U808 ( .A(reg_in_plain_text[72]), .Y(reg_in_n1010) );
  INVX1 reg_in_U807 ( .A(reg_in_plain_text[80]), .Y(reg_in_n1011) );
  INVX1 reg_in_U806 ( .A(reg_in_plain_text[88]), .Y(reg_in_n1012) );
  INVX1 reg_in_U805 ( .A(reg_in_plain_text[96]), .Y(reg_in_n1013) );
  INVX1 reg_in_U804 ( .A(reg_in_plain_text[104]), .Y(reg_in_n1014) );
  INVX1 reg_in_U803 ( .A(reg_in_plain_text[112]), .Y(reg_in_n1015) );
  INVX1 reg_in_U802 ( .A(reg_in_plain_text[120]), .Y(reg_in_n1016) );
  INVX1 reg_in_U801 ( .A(reg_in_plain_text[128]), .Y(reg_in_n1017) );
  INVX1 reg_in_U800 ( .A(reg_in_plain_text[136]), .Y(reg_in_n1018) );
  INVX1 reg_in_U799 ( .A(reg_in_plain_text[144]), .Y(reg_in_n1019) );
  INVX1 reg_in_U798 ( .A(reg_in_plain_text[152]), .Y(reg_in_n1020) );
  INVX1 reg_in_U797 ( .A(reg_in_plain_text[160]), .Y(reg_in_n1021) );
  INVX1 reg_in_U796 ( .A(reg_in_plain_text[168]), .Y(reg_in_n1022) );
  INVX1 reg_in_U795 ( .A(reg_in_plain_text[176]), .Y(reg_in_n1023) );
  INVX1 reg_in_U794 ( .A(reg_in_plain_text[184]), .Y(reg_in_n1024) );
  INVX1 reg_in_U793 ( .A(reg_in_plain_text[192]), .Y(reg_in_n1025) );
  INVX1 reg_in_U792 ( .A(reg_in_plain_text[200]), .Y(reg_in_n1026) );
  INVX1 reg_in_U791 ( .A(reg_in_plain_text[208]), .Y(reg_in_n1027) );
  INVX1 reg_in_U790 ( .A(reg_in_plain_text[216]), .Y(reg_in_n1028) );
  INVX1 reg_in_U789 ( .A(reg_in_plain_text[224]), .Y(reg_in_n1029) );
  INVX1 reg_in_U788 ( .A(reg_in_plain_text[232]), .Y(reg_in_n1030) );
  INVX1 reg_in_U787 ( .A(reg_in_plain_text[240]), .Y(reg_in_n1031) );
  INVX1 reg_in_U786 ( .A(reg_in_plain_text[7]), .Y(reg_in_n777) );
  INVX1 reg_in_U785 ( .A(reg_in_plain_text[6]), .Y(reg_in_n809) );
  INVX1 reg_in_U784 ( .A(reg_in_plain_text[5]), .Y(reg_in_n841) );
  INVX1 reg_in_U783 ( .A(reg_in_plain_text[4]), .Y(reg_in_n873) );
  INVX1 reg_in_U782 ( .A(reg_in_plain_text[3]), .Y(reg_in_n905) );
  INVX1 reg_in_U781 ( .A(reg_in_plain_text[2]), .Y(reg_in_n937) );
  INVX1 reg_in_U780 ( .A(reg_in_plain_text[1]), .Y(reg_in_n969) );
  INVX1 reg_in_U779 ( .A(reg_in_plain_text[0]), .Y(reg_in_n1001) );
  OAI2BB2X1 reg_in_U778 ( .B0(reg_in_n223), .B1(reg_in_n808), .A0N(Din[255]), 
        .A1N(reg_in_n251), .Y(reg_in_n515) );
  OAI2BB2X1 reg_in_U777 ( .B0(reg_in_n220), .B1(reg_in_n840), .A0N(Din[254]), 
        .A1N(reg_in_n250), .Y(reg_in_n514) );
  OAI2BB2X1 reg_in_U776 ( .B0(reg_in_n251), .B1(reg_in_n872), .A0N(Din[253]), 
        .A1N(reg_in_n240), .Y(reg_in_n513) );
  OAI2BB2X1 reg_in_U775 ( .B0(reg_in_n250), .B1(reg_in_n904), .A0N(Din[252]), 
        .A1N(reg_in_n240), .Y(reg_in_n512) );
  OAI2BB2X1 reg_in_U774 ( .B0(reg_in_n233), .B1(reg_in_n936), .A0N(Din[251]), 
        .A1N(reg_in_n240), .Y(reg_in_n511) );
  OAI2BB2X1 reg_in_U773 ( .B0(reg_in_n233), .B1(reg_in_n968), .A0N(Din[250]), 
        .A1N(reg_in_n240), .Y(reg_in_n510) );
  OAI2BB2X1 reg_in_U772 ( .B0(reg_in_n233), .B1(reg_in_n1000), .A0N(Din[249]), 
        .A1N(reg_in_n241), .Y(reg_in_n509) );
  OAI2BB2X1 reg_in_U771 ( .B0(reg_in_n233), .B1(reg_in_n1032), .A0N(Din[248]), 
        .A1N(reg_in_n242), .Y(reg_in_n508) );
  OAI2BB2X1 reg_in_U770 ( .B0(reg_in_n233), .B1(reg_in_n807), .A0N(Din[247]), 
        .A1N(reg_in_n241), .Y(reg_in_n507) );
  OAI2BB2X1 reg_in_U769 ( .B0(reg_in_n233), .B1(reg_in_n839), .A0N(Din[246]), 
        .A1N(reg_in_n241), .Y(reg_in_n506) );
  OAI2BB2X1 reg_in_U768 ( .B0(reg_in_n233), .B1(reg_in_n871), .A0N(Din[245]), 
        .A1N(reg_in_n242), .Y(reg_in_n505) );
  OAI2BB2X1 reg_in_U767 ( .B0(reg_in_n233), .B1(reg_in_n903), .A0N(Din[244]), 
        .A1N(reg_in_n242), .Y(reg_in_n504) );
  OAI2BB2X1 reg_in_U766 ( .B0(reg_in_n233), .B1(reg_in_n935), .A0N(Din[243]), 
        .A1N(reg_in_n242), .Y(reg_in_n503) );
  OAI2BB2X1 reg_in_U765 ( .B0(reg_in_n233), .B1(reg_in_n967), .A0N(Din[242]), 
        .A1N(reg_in_n243), .Y(reg_in_n502) );
  OAI2BB2X1 reg_in_U764 ( .B0(reg_in_n233), .B1(reg_in_n999), .A0N(Din[241]), 
        .A1N(reg_in_n243), .Y(reg_in_n501) );
  OAI2BB2X1 reg_in_U763 ( .B0(reg_in_n233), .B1(reg_in_n1031), .A0N(Din[240]), 
        .A1N(reg_in_n243), .Y(reg_in_n500) );
  OAI2BB2X1 reg_in_U762 ( .B0(reg_in_n232), .B1(reg_in_n806), .A0N(Din[239]), 
        .A1N(reg_in_n243), .Y(reg_in_n499) );
  OAI2BB2X1 reg_in_U761 ( .B0(reg_in_n232), .B1(reg_in_n838), .A0N(Din[238]), 
        .A1N(reg_in_n244), .Y(reg_in_n498) );
  OAI2BB2X1 reg_in_U760 ( .B0(reg_in_n232), .B1(reg_in_n870), .A0N(Din[237]), 
        .A1N(reg_in_n244), .Y(reg_in_n497) );
  OAI2BB2X1 reg_in_U759 ( .B0(reg_in_n232), .B1(reg_in_n902), .A0N(Din[236]), 
        .A1N(reg_in_n244), .Y(reg_in_n496) );
  OAI2BB2X1 reg_in_U758 ( .B0(reg_in_n232), .B1(reg_in_n934), .A0N(Din[235]), 
        .A1N(reg_in_n245), .Y(reg_in_n495) );
  OAI2BB2X1 reg_in_U757 ( .B0(reg_in_n232), .B1(reg_in_n966), .A0N(Din[234]), 
        .A1N(reg_in_n245), .Y(reg_in_n494) );
  OAI2BB2X1 reg_in_U756 ( .B0(reg_in_n232), .B1(reg_in_n998), .A0N(Din[233]), 
        .A1N(reg_in_n245), .Y(reg_in_n493) );
  OAI2BB2X1 reg_in_U755 ( .B0(reg_in_n232), .B1(reg_in_n1030), .A0N(Din[232]), 
        .A1N(reg_in_n245), .Y(reg_in_n492) );
  OAI2BB2X1 reg_in_U754 ( .B0(reg_in_n232), .B1(reg_in_n805), .A0N(Din[231]), 
        .A1N(reg_in_n245), .Y(reg_in_n491) );
  OAI2BB2X1 reg_in_U753 ( .B0(reg_in_n232), .B1(reg_in_n837), .A0N(Din[230]), 
        .A1N(reg_in_n245), .Y(reg_in_n490) );
  OAI2BB2X1 reg_in_U752 ( .B0(reg_in_n232), .B1(reg_in_n869), .A0N(Din[229]), 
        .A1N(reg_in_n244), .Y(reg_in_n489) );
  OAI2BB2X1 reg_in_U751 ( .B0(reg_in_n232), .B1(reg_in_n901), .A0N(Din[228]), 
        .A1N(reg_in_n244), .Y(reg_in_n488) );
  OAI2BB2X1 reg_in_U750 ( .B0(reg_in_n231), .B1(reg_in_n933), .A0N(Din[227]), 
        .A1N(reg_in_n244), .Y(reg_in_n487) );
  OAI2BB2X1 reg_in_U749 ( .B0(reg_in_n231), .B1(reg_in_n965), .A0N(Din[226]), 
        .A1N(reg_in_n244), .Y(reg_in_n486) );
  OAI2BB2X1 reg_in_U748 ( .B0(reg_in_n231), .B1(reg_in_n997), .A0N(Din[225]), 
        .A1N(reg_in_n244), .Y(reg_in_n485) );
  OAI2BB2X1 reg_in_U747 ( .B0(reg_in_n231), .B1(reg_in_n1029), .A0N(Din[224]), 
        .A1N(reg_in_n244), .Y(reg_in_n484) );
  OAI2BB2X1 reg_in_U746 ( .B0(reg_in_n231), .B1(reg_in_n804), .A0N(Din[223]), 
        .A1N(reg_in_n244), .Y(reg_in_n483) );
  OAI2BB2X1 reg_in_U745 ( .B0(reg_in_n231), .B1(reg_in_n836), .A0N(Din[222]), 
        .A1N(reg_in_n244), .Y(reg_in_n482) );
  OAI2BB2X1 reg_in_U744 ( .B0(reg_in_n231), .B1(reg_in_n868), .A0N(Din[221]), 
        .A1N(reg_in_n244), .Y(reg_in_n481) );
  OAI2BB2X1 reg_in_U743 ( .B0(reg_in_n231), .B1(reg_in_n900), .A0N(Din[220]), 
        .A1N(reg_in_n243), .Y(reg_in_n480) );
  OAI2BB2X1 reg_in_U742 ( .B0(reg_in_n231), .B1(reg_in_n932), .A0N(Din[219]), 
        .A1N(reg_in_n243), .Y(reg_in_n479) );
  OAI2BB2X1 reg_in_U741 ( .B0(reg_in_n231), .B1(reg_in_n964), .A0N(Din[218]), 
        .A1N(reg_in_n243), .Y(reg_in_n478) );
  OAI2BB2X1 reg_in_U740 ( .B0(reg_in_n231), .B1(reg_in_n996), .A0N(Din[217]), 
        .A1N(reg_in_n243), .Y(reg_in_n477) );
  OAI2BB2X1 reg_in_U739 ( .B0(reg_in_n231), .B1(reg_in_n1028), .A0N(Din[216]), 
        .A1N(reg_in_n243), .Y(reg_in_n476) );
  OAI2BB2X1 reg_in_U738 ( .B0(reg_in_n230), .B1(reg_in_n803), .A0N(Din[215]), 
        .A1N(reg_in_n243), .Y(reg_in_n475) );
  OAI2BB2X1 reg_in_U737 ( .B0(reg_in_n230), .B1(reg_in_n835), .A0N(Din[214]), 
        .A1N(reg_in_n243), .Y(reg_in_n474) );
  OAI2BB2X1 reg_in_U736 ( .B0(reg_in_n230), .B1(reg_in_n867), .A0N(Din[213]), 
        .A1N(reg_in_n243), .Y(reg_in_n473) );
  OAI2BB2X1 reg_in_U735 ( .B0(reg_in_n230), .B1(reg_in_n899), .A0N(Din[212]), 
        .A1N(reg_in_n242), .Y(reg_in_n472) );
  OAI2BB2X1 reg_in_U734 ( .B0(reg_in_n230), .B1(reg_in_n931), .A0N(Din[211]), 
        .A1N(reg_in_n242), .Y(reg_in_n471) );
  OAI2BB2X1 reg_in_U733 ( .B0(reg_in_n230), .B1(reg_in_n963), .A0N(Din[210]), 
        .A1N(reg_in_n242), .Y(reg_in_n470) );
  OAI2BB2X1 reg_in_U732 ( .B0(reg_in_n230), .B1(reg_in_n995), .A0N(Din[209]), 
        .A1N(reg_in_n242), .Y(reg_in_n469) );
  OAI2BB2X1 reg_in_U731 ( .B0(reg_in_n230), .B1(reg_in_n1027), .A0N(Din[208]), 
        .A1N(reg_in_n242), .Y(reg_in_n468) );
  OAI2BB2X1 reg_in_U730 ( .B0(reg_in_n230), .B1(reg_in_n802), .A0N(Din[207]), 
        .A1N(reg_in_n242), .Y(reg_in_n467) );
  OAI2BB2X1 reg_in_U729 ( .B0(reg_in_n230), .B1(reg_in_n834), .A0N(Din[206]), 
        .A1N(reg_in_n242), .Y(reg_in_n466) );
  OAI2BB2X1 reg_in_U728 ( .B0(reg_in_n230), .B1(reg_in_n866), .A0N(Din[205]), 
        .A1N(reg_in_n241), .Y(reg_in_n465) );
  OAI2BB2X1 reg_in_U727 ( .B0(reg_in_n230), .B1(reg_in_n898), .A0N(Din[204]), 
        .A1N(reg_in_n241), .Y(reg_in_n464) );
  OAI2BB2X1 reg_in_U726 ( .B0(reg_in_n229), .B1(reg_in_n930), .A0N(Din[203]), 
        .A1N(reg_in_n241), .Y(reg_in_n463) );
  OAI2BB2X1 reg_in_U725 ( .B0(reg_in_n229), .B1(reg_in_n962), .A0N(Din[202]), 
        .A1N(reg_in_n241), .Y(reg_in_n462) );
  OAI2BB2X1 reg_in_U724 ( .B0(reg_in_n229), .B1(reg_in_n994), .A0N(Din[201]), 
        .A1N(reg_in_n241), .Y(reg_in_n461) );
  OAI2BB2X1 reg_in_U723 ( .B0(reg_in_n229), .B1(reg_in_n1026), .A0N(Din[200]), 
        .A1N(reg_in_n241), .Y(reg_in_n460) );
  OAI2BB2X1 reg_in_U722 ( .B0(reg_in_n229), .B1(reg_in_n801), .A0N(Din[199]), 
        .A1N(reg_in_n240), .Y(reg_in_n459) );
  OAI2BB2X1 reg_in_U721 ( .B0(reg_in_n229), .B1(reg_in_n833), .A0N(Din[198]), 
        .A1N(reg_in_n240), .Y(reg_in_n458) );
  OAI2BB2X1 reg_in_U720 ( .B0(reg_in_n229), .B1(reg_in_n865), .A0N(Din[197]), 
        .A1N(reg_in_n241), .Y(reg_in_n457) );
  OAI2BB2X1 reg_in_U719 ( .B0(reg_in_n229), .B1(reg_in_n897), .A0N(Din[196]), 
        .A1N(reg_in_n241), .Y(reg_in_n456) );
  OAI2BB2X1 reg_in_U718 ( .B0(reg_in_n229), .B1(reg_in_n929), .A0N(Din[195]), 
        .A1N(reg_in_n240), .Y(reg_in_n455) );
  OAI2BB2X1 reg_in_U717 ( .B0(reg_in_n229), .B1(reg_in_n961), .A0N(Din[194]), 
        .A1N(reg_in_n240), .Y(reg_in_n454) );
  OAI2BB2X1 reg_in_U716 ( .B0(reg_in_n229), .B1(reg_in_n993), .A0N(Din[193]), 
        .A1N(reg_in_n240), .Y(reg_in_n453) );
  OAI2BB2X1 reg_in_U715 ( .B0(reg_in_n229), .B1(reg_in_n1025), .A0N(Din[192]), 
        .A1N(reg_in_n241), .Y(reg_in_n452) );
  OAI2BB2X1 reg_in_U714 ( .B0(reg_in_n228), .B1(reg_in_n800), .A0N(Din[191]), 
        .A1N(reg_in_n249), .Y(reg_in_n451) );
  OAI2BB2X1 reg_in_U713 ( .B0(reg_in_n228), .B1(reg_in_n832), .A0N(Din[190]), 
        .A1N(reg_in_n240), .Y(reg_in_n450) );
  OAI2BB2X1 reg_in_U712 ( .B0(reg_in_n228), .B1(reg_in_n864), .A0N(Din[189]), 
        .A1N(reg_in_n240), .Y(reg_in_n449) );
  OAI2BB2X1 reg_in_U711 ( .B0(reg_in_n228), .B1(reg_in_n896), .A0N(Din[188]), 
        .A1N(reg_in_n248), .Y(reg_in_n448) );
  OAI2BB2X1 reg_in_U710 ( .B0(reg_in_n228), .B1(reg_in_n928), .A0N(Din[187]), 
        .A1N(reg_in_n241), .Y(reg_in_n447) );
  OAI2BB2X1 reg_in_U709 ( .B0(reg_in_n228), .B1(reg_in_n960), .A0N(Din[186]), 
        .A1N(reg_in_n240), .Y(reg_in_n446) );
  OAI2BB2X1 reg_in_U708 ( .B0(reg_in_n228), .B1(reg_in_n992), .A0N(Din[185]), 
        .A1N(reg_in_n240), .Y(reg_in_n445) );
  OAI2BB2X1 reg_in_U707 ( .B0(reg_in_n228), .B1(reg_in_n1024), .A0N(Din[184]), 
        .A1N(reg_in_n241), .Y(reg_in_n444) );
  OAI2BB2X1 reg_in_U706 ( .B0(reg_in_n228), .B1(reg_in_n799), .A0N(Din[183]), 
        .A1N(reg_in_n252), .Y(reg_in_n443) );
  OAI2BB2X1 reg_in_U705 ( .B0(reg_in_n228), .B1(reg_in_n831), .A0N(Din[182]), 
        .A1N(reg_in_n253), .Y(reg_in_n442) );
  OAI2BB2X1 reg_in_U704 ( .B0(reg_in_n228), .B1(reg_in_n863), .A0N(Din[181]), 
        .A1N(reg_in_n253), .Y(reg_in_n441) );
  OAI2BB2X1 reg_in_U703 ( .B0(reg_in_n228), .B1(reg_in_n895), .A0N(Din[180]), 
        .A1N(reg_in_n253), .Y(reg_in_n440) );
  OAI2BB2X1 reg_in_U702 ( .B0(reg_in_n227), .B1(reg_in_n927), .A0N(Din[179]), 
        .A1N(reg_in_n253), .Y(reg_in_n439) );
  OAI2BB2X1 reg_in_U701 ( .B0(reg_in_n227), .B1(reg_in_n959), .A0N(Din[178]), 
        .A1N(reg_in_n253), .Y(reg_in_n438) );
  OAI2BB2X1 reg_in_U700 ( .B0(reg_in_n227), .B1(reg_in_n991), .A0N(Din[177]), 
        .A1N(reg_in_n253), .Y(reg_in_n437) );
  OAI2BB2X1 reg_in_U699 ( .B0(reg_in_n227), .B1(reg_in_n1023), .A0N(Din[176]), 
        .A1N(reg_in_n253), .Y(reg_in_n436) );
  OAI2BB2X1 reg_in_U698 ( .B0(reg_in_n227), .B1(reg_in_n798), .A0N(Din[175]), 
        .A1N(reg_in_n252), .Y(reg_in_n435) );
  OAI2BB2X1 reg_in_U697 ( .B0(reg_in_n227), .B1(reg_in_n830), .A0N(Din[174]), 
        .A1N(reg_in_n252), .Y(reg_in_n434) );
  OAI2BB2X1 reg_in_U696 ( .B0(reg_in_n227), .B1(reg_in_n862), .A0N(Din[173]), 
        .A1N(reg_in_n252), .Y(reg_in_n433) );
  OAI2BB2X1 reg_in_U695 ( .B0(reg_in_n227), .B1(reg_in_n894), .A0N(Din[172]), 
        .A1N(reg_in_n252), .Y(reg_in_n432) );
  OAI2BB2X1 reg_in_U694 ( .B0(reg_in_n227), .B1(reg_in_n926), .A0N(Din[171]), 
        .A1N(reg_in_n252), .Y(reg_in_n431) );
  OAI2BB2X1 reg_in_U693 ( .B0(reg_in_n227), .B1(reg_in_n958), .A0N(Din[170]), 
        .A1N(reg_in_n252), .Y(reg_in_n430) );
  OAI2BB2X1 reg_in_U692 ( .B0(reg_in_n227), .B1(reg_in_n990), .A0N(Din[169]), 
        .A1N(reg_in_n252), .Y(reg_in_n429) );
  OAI2BB2X1 reg_in_U691 ( .B0(reg_in_n226), .B1(reg_in_n1022), .A0N(Din[168]), 
        .A1N(reg_in_n252), .Y(reg_in_n428) );
  OAI2BB2X1 reg_in_U690 ( .B0(reg_in_n226), .B1(reg_in_n797), .A0N(Din[167]), 
        .A1N(reg_in_n252), .Y(reg_in_n427) );
  OAI2BB2X1 reg_in_U689 ( .B0(reg_in_n226), .B1(reg_in_n829), .A0N(Din[166]), 
        .A1N(reg_in_n252), .Y(reg_in_n426) );
  OAI2BB2X1 reg_in_U688 ( .B0(reg_in_n226), .B1(reg_in_n861), .A0N(Din[165]), 
        .A1N(reg_in_n252), .Y(reg_in_n425) );
  OAI2BB2X1 reg_in_U687 ( .B0(reg_in_n226), .B1(reg_in_n893), .A0N(Din[164]), 
        .A1N(reg_in_n252), .Y(reg_in_n424) );
  OAI2BB2X1 reg_in_U686 ( .B0(reg_in_n226), .B1(reg_in_n925), .A0N(Din[163]), 
        .A1N(reg_in_n251), .Y(reg_in_n423) );
  OAI2BB2X1 reg_in_U685 ( .B0(reg_in_n226), .B1(reg_in_n957), .A0N(Din[162]), 
        .A1N(reg_in_n251), .Y(reg_in_n422) );
  OAI2BB2X1 reg_in_U684 ( .B0(reg_in_n226), .B1(reg_in_n989), .A0N(Din[161]), 
        .A1N(reg_in_n251), .Y(reg_in_n421) );
  OAI2BB2X1 reg_in_U683 ( .B0(reg_in_n226), .B1(reg_in_n1021), .A0N(Din[160]), 
        .A1N(reg_in_n251), .Y(reg_in_n420) );
  OAI2BB2X1 reg_in_U682 ( .B0(reg_in_n226), .B1(reg_in_n796), .A0N(Din[159]), 
        .A1N(reg_in_n251), .Y(reg_in_n419) );
  OAI2BB2X1 reg_in_U681 ( .B0(reg_in_n226), .B1(reg_in_n828), .A0N(Din[158]), 
        .A1N(reg_in_n251), .Y(reg_in_n418) );
  OAI2BB2X1 reg_in_U680 ( .B0(reg_in_n226), .B1(reg_in_n860), .A0N(Din[157]), 
        .A1N(reg_in_n251), .Y(reg_in_n417) );
  OAI2BB2X1 reg_in_U679 ( .B0(reg_in_n225), .B1(reg_in_n892), .A0N(Din[156]), 
        .A1N(reg_in_n251), .Y(reg_in_n416) );
  OAI2BB2X1 reg_in_U678 ( .B0(reg_in_n225), .B1(reg_in_n924), .A0N(Din[155]), 
        .A1N(reg_in_n251), .Y(reg_in_n415) );
  OAI2BB2X1 reg_in_U677 ( .B0(reg_in_n225), .B1(reg_in_n956), .A0N(Din[154]), 
        .A1N(reg_in_n251), .Y(reg_in_n414) );
  OAI2BB2X1 reg_in_U676 ( .B0(reg_in_n225), .B1(reg_in_n988), .A0N(Din[153]), 
        .A1N(reg_in_n251), .Y(reg_in_n413) );
  OAI2BB2X1 reg_in_U675 ( .B0(reg_in_n225), .B1(reg_in_n1020), .A0N(Din[152]), 
        .A1N(reg_in_n251), .Y(reg_in_n412) );
  OAI2BB2X1 reg_in_U674 ( .B0(reg_in_n225), .B1(reg_in_n795), .A0N(Din[151]), 
        .A1N(reg_in_n250), .Y(reg_in_n411) );
  OAI2BB2X1 reg_in_U673 ( .B0(reg_in_n225), .B1(reg_in_n827), .A0N(Din[150]), 
        .A1N(reg_in_n250), .Y(reg_in_n410) );
  OAI2BB2X1 reg_in_U672 ( .B0(reg_in_n225), .B1(reg_in_n859), .A0N(Din[149]), 
        .A1N(reg_in_n250), .Y(reg_in_n409) );
  OAI2BB2X1 reg_in_U671 ( .B0(reg_in_n225), .B1(reg_in_n891), .A0N(Din[148]), 
        .A1N(reg_in_n250), .Y(reg_in_n408) );
  OAI2BB2X1 reg_in_U670 ( .B0(reg_in_n225), .B1(reg_in_n923), .A0N(Din[147]), 
        .A1N(reg_in_n250), .Y(reg_in_n407) );
  OAI2BB2X1 reg_in_U669 ( .B0(reg_in_n225), .B1(reg_in_n955), .A0N(Din[146]), 
        .A1N(reg_in_n250), .Y(reg_in_n406) );
  OAI2BB2X1 reg_in_U668 ( .B0(reg_in_n225), .B1(reg_in_n987), .A0N(Din[145]), 
        .A1N(reg_in_n250), .Y(reg_in_n405) );
  OAI2BB2X1 reg_in_U667 ( .B0(reg_in_n224), .B1(reg_in_n1019), .A0N(Din[144]), 
        .A1N(reg_in_n250), .Y(reg_in_n404) );
  OAI2BB2X1 reg_in_U666 ( .B0(reg_in_n224), .B1(reg_in_n794), .A0N(Din[143]), 
        .A1N(reg_in_n250), .Y(reg_in_n403) );
  OAI2BB2X1 reg_in_U665 ( .B0(reg_in_n224), .B1(reg_in_n826), .A0N(Din[142]), 
        .A1N(reg_in_n250), .Y(reg_in_n402) );
  OAI2BB2X1 reg_in_U664 ( .B0(reg_in_n224), .B1(reg_in_n858), .A0N(Din[141]), 
        .A1N(reg_in_n250), .Y(reg_in_n401) );
  OAI2BB2X1 reg_in_U663 ( .B0(reg_in_n224), .B1(reg_in_n890), .A0N(Din[140]), 
        .A1N(reg_in_n250), .Y(reg_in_n400) );
  OAI2BB2X1 reg_in_U662 ( .B0(reg_in_n224), .B1(reg_in_n922), .A0N(Din[139]), 
        .A1N(reg_in_n249), .Y(reg_in_n399) );
  OAI2BB2X1 reg_in_U661 ( .B0(reg_in_n224), .B1(reg_in_n954), .A0N(Din[138]), 
        .A1N(reg_in_n249), .Y(reg_in_n398) );
  OAI2BB2X1 reg_in_U660 ( .B0(reg_in_n224), .B1(reg_in_n986), .A0N(Din[137]), 
        .A1N(reg_in_n249), .Y(reg_in_n397) );
  OAI2BB2X1 reg_in_U659 ( .B0(reg_in_n224), .B1(reg_in_n1018), .A0N(Din[136]), 
        .A1N(reg_in_n249), .Y(reg_in_n396) );
  OAI2BB2X1 reg_in_U658 ( .B0(reg_in_n224), .B1(reg_in_n793), .A0N(Din[135]), 
        .A1N(reg_in_n249), .Y(reg_in_n395) );
  OAI2BB2X1 reg_in_U657 ( .B0(reg_in_n224), .B1(reg_in_n825), .A0N(Din[134]), 
        .A1N(reg_in_n249), .Y(reg_in_n394) );
  OAI2BB2X1 reg_in_U656 ( .B0(reg_in_n224), .B1(reg_in_n857), .A0N(Din[133]), 
        .A1N(reg_in_n249), .Y(reg_in_n393) );
  OAI2BB2X1 reg_in_U655 ( .B0(reg_in_n223), .B1(reg_in_n889), .A0N(Din[132]), 
        .A1N(reg_in_n249), .Y(reg_in_n392) );
  OAI2BB2X1 reg_in_U654 ( .B0(reg_in_n223), .B1(reg_in_n921), .A0N(Din[131]), 
        .A1N(reg_in_n249), .Y(reg_in_n391) );
  OAI2BB2X1 reg_in_U653 ( .B0(reg_in_n223), .B1(reg_in_n953), .A0N(Din[130]), 
        .A1N(reg_in_n249), .Y(reg_in_n390) );
  OAI2BB2X1 reg_in_U652 ( .B0(reg_in_n223), .B1(reg_in_n985), .A0N(Din[129]), 
        .A1N(reg_in_n249), .Y(reg_in_n389) );
  OAI2BB2X1 reg_in_U651 ( .B0(reg_in_n223), .B1(reg_in_n1017), .A0N(Din[128]), 
        .A1N(reg_in_n248), .Y(reg_in_n388) );
  OAI2BB2X1 reg_in_U650 ( .B0(reg_in_n240), .B1(reg_in_n792), .A0N(Din[127]), 
        .A1N(reg_in_n248), .Y(reg_in_n387) );
  OAI2BB2X1 reg_in_U649 ( .B0(reg_in_n223), .B1(reg_in_n824), .A0N(Din[126]), 
        .A1N(reg_in_n248), .Y(reg_in_n386) );
  OAI2BB2X1 reg_in_U648 ( .B0(reg_in_n223), .B1(reg_in_n856), .A0N(Din[125]), 
        .A1N(reg_in_n248), .Y(reg_in_n385) );
  OAI2BB2X1 reg_in_U647 ( .B0(reg_in_n223), .B1(reg_in_n888), .A0N(Din[124]), 
        .A1N(reg_in_n248), .Y(reg_in_n384) );
  OAI2BB2X1 reg_in_U646 ( .B0(reg_in_n223), .B1(reg_in_n920), .A0N(Din[123]), 
        .A1N(reg_in_n248), .Y(reg_in_n383) );
  OAI2BB2X1 reg_in_U645 ( .B0(reg_in_n223), .B1(reg_in_n952), .A0N(Din[122]), 
        .A1N(reg_in_n248), .Y(reg_in_n382) );
  OAI2BB2X1 reg_in_U644 ( .B0(reg_in_n223), .B1(reg_in_n984), .A0N(Din[121]), 
        .A1N(reg_in_n248), .Y(reg_in_n381) );
  OAI2BB2X1 reg_in_U643 ( .B0(reg_in_n222), .B1(reg_in_n1016), .A0N(Din[120]), 
        .A1N(reg_in_n248), .Y(reg_in_n380) );
  OAI2BB2X1 reg_in_U642 ( .B0(reg_in_n222), .B1(reg_in_n791), .A0N(Din[119]), 
        .A1N(reg_in_n248), .Y(reg_in_n379) );
  OAI2BB2X1 reg_in_U641 ( .B0(reg_in_n222), .B1(reg_in_n823), .A0N(Din[118]), 
        .A1N(reg_in_n248), .Y(reg_in_n378) );
  OAI2BB2X1 reg_in_U640 ( .B0(reg_in_n222), .B1(reg_in_n855), .A0N(Din[117]), 
        .A1N(reg_in_n248), .Y(reg_in_n377) );
  OAI2BB2X1 reg_in_U639 ( .B0(reg_in_n222), .B1(reg_in_n887), .A0N(Din[116]), 
        .A1N(reg_in_n247), .Y(reg_in_n376) );
  OAI2BB2X1 reg_in_U638 ( .B0(reg_in_n222), .B1(reg_in_n919), .A0N(Din[115]), 
        .A1N(reg_in_n247), .Y(reg_in_n375) );
  OAI2BB2X1 reg_in_U637 ( .B0(reg_in_n222), .B1(reg_in_n951), .A0N(Din[114]), 
        .A1N(reg_in_n247), .Y(reg_in_n374) );
  OAI2BB2X1 reg_in_U636 ( .B0(reg_in_n222), .B1(reg_in_n983), .A0N(Din[113]), 
        .A1N(reg_in_n247), .Y(reg_in_n373) );
  OAI2BB2X1 reg_in_U635 ( .B0(reg_in_n222), .B1(reg_in_n1015), .A0N(Din[112]), 
        .A1N(reg_in_n247), .Y(reg_in_n372) );
  OAI2BB2X1 reg_in_U634 ( .B0(reg_in_n222), .B1(reg_in_n790), .A0N(Din[111]), 
        .A1N(reg_in_n247), .Y(reg_in_n371) );
  OAI2BB2X1 reg_in_U633 ( .B0(reg_in_n222), .B1(reg_in_n822), .A0N(Din[110]), 
        .A1N(reg_in_n247), .Y(reg_in_n370) );
  OAI2BB2X1 reg_in_U632 ( .B0(reg_in_n222), .B1(reg_in_n854), .A0N(Din[109]), 
        .A1N(reg_in_n247), .Y(reg_in_n369) );
  OAI2BB2X1 reg_in_U631 ( .B0(reg_in_n221), .B1(reg_in_n886), .A0N(Din[108]), 
        .A1N(reg_in_n247), .Y(reg_in_n368) );
  OAI2BB2X1 reg_in_U630 ( .B0(reg_in_n221), .B1(reg_in_n918), .A0N(Din[107]), 
        .A1N(reg_in_n247), .Y(reg_in_n367) );
  OAI2BB2X1 reg_in_U629 ( .B0(reg_in_n221), .B1(reg_in_n950), .A0N(Din[106]), 
        .A1N(reg_in_n247), .Y(reg_in_n366) );
  OAI2BB2X1 reg_in_U628 ( .B0(reg_in_n221), .B1(reg_in_n982), .A0N(Din[105]), 
        .A1N(reg_in_n247), .Y(reg_in_n365) );
  OAI2BB2X1 reg_in_U627 ( .B0(reg_in_n221), .B1(reg_in_n1014), .A0N(Din[104]), 
        .A1N(reg_in_n246), .Y(reg_in_n364) );
  OAI2BB2X1 reg_in_U626 ( .B0(reg_in_n221), .B1(reg_in_n789), .A0N(Din[103]), 
        .A1N(reg_in_n246), .Y(reg_in_n363) );
  OAI2BB2X1 reg_in_U625 ( .B0(reg_in_n221), .B1(reg_in_n821), .A0N(Din[102]), 
        .A1N(reg_in_n246), .Y(reg_in_n362) );
  OAI2BB2X1 reg_in_U624 ( .B0(reg_in_n221), .B1(reg_in_n853), .A0N(Din[101]), 
        .A1N(reg_in_n246), .Y(reg_in_n361) );
  OAI2BB2X1 reg_in_U623 ( .B0(reg_in_n221), .B1(reg_in_n885), .A0N(Din[100]), 
        .A1N(reg_in_n246), .Y(reg_in_n360) );
  OAI2BB2X1 reg_in_U622 ( .B0(reg_in_n221), .B1(reg_in_n917), .A0N(Din[99]), 
        .A1N(reg_in_n246), .Y(reg_in_n359) );
  OAI2BB2X1 reg_in_U621 ( .B0(reg_in_n221), .B1(reg_in_n949), .A0N(Din[98]), 
        .A1N(reg_in_n246), .Y(reg_in_n358) );
  OAI2BB2X1 reg_in_U620 ( .B0(reg_in_n221), .B1(reg_in_n981), .A0N(Din[97]), 
        .A1N(reg_in_n246), .Y(reg_in_n357) );
  OAI2BB2X1 reg_in_U619 ( .B0(reg_in_n220), .B1(reg_in_n1013), .A0N(Din[96]), 
        .A1N(reg_in_n246), .Y(reg_in_n356) );
  OAI2BB2X1 reg_in_U618 ( .B0(reg_in_n220), .B1(reg_in_n788), .A0N(Din[95]), 
        .A1N(reg_in_n246), .Y(reg_in_n355) );
  OAI2BB2X1 reg_in_U617 ( .B0(reg_in_n220), .B1(reg_in_n820), .A0N(Din[94]), 
        .A1N(reg_in_n246), .Y(reg_in_n354) );
  OAI2BB2X1 reg_in_U616 ( .B0(reg_in_n220), .B1(reg_in_n852), .A0N(Din[93]), 
        .A1N(reg_in_n246), .Y(reg_in_n353) );
  OAI2BB2X1 reg_in_U615 ( .B0(reg_in_n220), .B1(reg_in_n884), .A0N(Din[92]), 
        .A1N(reg_in_n245), .Y(reg_in_n352) );
  OAI2BB2X1 reg_in_U614 ( .B0(reg_in_n220), .B1(reg_in_n916), .A0N(Din[91]), 
        .A1N(reg_in_n245), .Y(reg_in_n351) );
  OAI2BB2X1 reg_in_U613 ( .B0(reg_in_n220), .B1(reg_in_n948), .A0N(Din[90]), 
        .A1N(reg_in_n245), .Y(reg_in_n350) );
  OAI2BB2X1 reg_in_U612 ( .B0(reg_in_n220), .B1(reg_in_n980), .A0N(Din[89]), 
        .A1N(reg_in_n245), .Y(reg_in_n349) );
  OAI2BB2X1 reg_in_U611 ( .B0(reg_in_n220), .B1(reg_in_n1012), .A0N(Din[88]), 
        .A1N(reg_in_n245), .Y(reg_in_n348) );
  OAI2BB2X1 reg_in_U610 ( .B0(reg_in_n220), .B1(reg_in_n787), .A0N(Din[87]), 
        .A1N(reg_in_n245), .Y(reg_in_n347) );
  OAI2BB2X1 reg_in_U609 ( .B0(reg_in_n220), .B1(reg_in_n819), .A0N(Din[86]), 
        .A1N(reg_in_n249), .Y(reg_in_n346) );
  OAI2BB2X1 reg_in_U608 ( .B0(reg_in_n227), .B1(reg_in_n851), .A0N(Din[85]), 
        .A1N(reg_in_n242), .Y(reg_in_n345) );
  OAI2BB2X1 reg_in_U607 ( .B0(reg_in_n238), .B1(reg_in_n883), .A0N(Din[84]), 
        .A1N(reg_in_n245), .Y(reg_in_n344) );
  OAI2BB2X1 reg_in_U606 ( .B0(reg_in_n238), .B1(reg_in_n915), .A0N(Din[83]), 
        .A1N(reg_in_n245), .Y(reg_in_n343) );
  OAI2BB2X1 reg_in_U605 ( .B0(reg_in_n239), .B1(reg_in_n947), .A0N(Din[82]), 
        .A1N(reg_in_n245), .Y(reg_in_n342) );
  OAI2BB2X1 reg_in_U604 ( .B0(reg_in_n239), .B1(reg_in_n979), .A0N(Din[81]), 
        .A1N(reg_in_n246), .Y(reg_in_n341) );
  OAI2BB2X1 reg_in_U603 ( .B0(reg_in_n239), .B1(reg_in_n1011), .A0N(Din[80]), 
        .A1N(reg_in_n246), .Y(reg_in_n340) );
  OAI2BB2X1 reg_in_U602 ( .B0(reg_in_n239), .B1(reg_in_n786), .A0N(Din[79]), 
        .A1N(reg_in_n246), .Y(reg_in_n339) );
  OAI2BB2X1 reg_in_U601 ( .B0(reg_in_n239), .B1(reg_in_n818), .A0N(Din[78]), 
        .A1N(reg_in_n246), .Y(reg_in_n338) );
  OAI2BB2X1 reg_in_U600 ( .B0(reg_in_n239), .B1(reg_in_n850), .A0N(Din[77]), 
        .A1N(reg_in_n246), .Y(reg_in_n337) );
  OAI2BB2X1 reg_in_U599 ( .B0(reg_in_n238), .B1(reg_in_n882), .A0N(Din[76]), 
        .A1N(reg_in_n246), .Y(reg_in_n336) );
  OAI2BB2X1 reg_in_U598 ( .B0(reg_in_n242), .B1(reg_in_n914), .A0N(Din[75]), 
        .A1N(reg_in_n247), .Y(reg_in_n335) );
  OAI2BB2X1 reg_in_U597 ( .B0(reg_in_n239), .B1(reg_in_n946), .A0N(Din[74]), 
        .A1N(reg_in_n247), .Y(reg_in_n334) );
  OAI2BB2X1 reg_in_U596 ( .B0(reg_in_n238), .B1(reg_in_n978), .A0N(Din[73]), 
        .A1N(reg_in_n247), .Y(reg_in_n333) );
  OAI2BB2X1 reg_in_U595 ( .B0(reg_in_n239), .B1(reg_in_n1010), .A0N(Din[72]), 
        .A1N(reg_in_n247), .Y(reg_in_n332) );
  OAI2BB2X1 reg_in_U594 ( .B0(reg_in_n238), .B1(reg_in_n785), .A0N(Din[71]), 
        .A1N(reg_in_n247), .Y(reg_in_n331) );
  OAI2BB2X1 reg_in_U593 ( .B0(reg_in_n238), .B1(reg_in_n817), .A0N(Din[70]), 
        .A1N(reg_in_n247), .Y(reg_in_n330) );
  OAI2BB2X1 reg_in_U592 ( .B0(reg_in_n237), .B1(reg_in_n849), .A0N(Din[69]), 
        .A1N(reg_in_n248), .Y(reg_in_n329) );
  OAI2BB2X1 reg_in_U591 ( .B0(reg_in_n237), .B1(reg_in_n881), .A0N(Din[68]), 
        .A1N(reg_in_n248), .Y(reg_in_n328) );
  OAI2BB2X1 reg_in_U590 ( .B0(reg_in_n237), .B1(reg_in_n913), .A0N(Din[67]), 
        .A1N(reg_in_n248), .Y(reg_in_n327) );
  OAI2BB2X1 reg_in_U589 ( .B0(reg_in_n237), .B1(reg_in_n945), .A0N(Din[66]), 
        .A1N(reg_in_n248), .Y(reg_in_n326) );
  OAI2BB2X1 reg_in_U588 ( .B0(reg_in_n237), .B1(reg_in_n977), .A0N(Din[65]), 
        .A1N(reg_in_n248), .Y(reg_in_n325) );
  OAI2BB2X1 reg_in_U587 ( .B0(reg_in_n237), .B1(reg_in_n1009), .A0N(Din[64]), 
        .A1N(reg_in_n248), .Y(reg_in_n324) );
  OAI2BB2X1 reg_in_U586 ( .B0(reg_in_n237), .B1(reg_in_n784), .A0N(Din[63]), 
        .A1N(reg_in_n249), .Y(reg_in_n323) );
  OAI2BB2X1 reg_in_U585 ( .B0(reg_in_n236), .B1(reg_in_n816), .A0N(Din[62]), 
        .A1N(reg_in_n249), .Y(reg_in_n322) );
  OAI2BB2X1 reg_in_U584 ( .B0(reg_in_n236), .B1(reg_in_n848), .A0N(Din[61]), 
        .A1N(reg_in_n249), .Y(reg_in_n321) );
  OAI2BB2X1 reg_in_U583 ( .B0(reg_in_n236), .B1(reg_in_n880), .A0N(Din[60]), 
        .A1N(reg_in_n249), .Y(reg_in_n320) );
  OAI2BB2X1 reg_in_U582 ( .B0(reg_in_n236), .B1(reg_in_n912), .A0N(Din[59]), 
        .A1N(reg_in_n249), .Y(reg_in_n319) );
  OAI2BB2X1 reg_in_U581 ( .B0(reg_in_n236), .B1(reg_in_n944), .A0N(Din[58]), 
        .A1N(reg_in_n249), .Y(reg_in_n318) );
  OAI2BB2X1 reg_in_U580 ( .B0(reg_in_n236), .B1(reg_in_n976), .A0N(Din[57]), 
        .A1N(reg_in_n250), .Y(reg_in_n317) );
  OAI2BB2X1 reg_in_U579 ( .B0(reg_in_n236), .B1(reg_in_n1008), .A0N(Din[56]), 
        .A1N(reg_in_n250), .Y(reg_in_n316) );
  OAI2BB2X1 reg_in_U578 ( .B0(reg_in_n235), .B1(reg_in_n783), .A0N(Din[55]), 
        .A1N(reg_in_n250), .Y(reg_in_n315) );
  OAI2BB2X1 reg_in_U577 ( .B0(reg_in_n235), .B1(reg_in_n815), .A0N(Din[54]), 
        .A1N(reg_in_n250), .Y(reg_in_n314) );
  OAI2BB2X1 reg_in_U576 ( .B0(reg_in_n235), .B1(reg_in_n847), .A0N(Din[53]), 
        .A1N(reg_in_n250), .Y(reg_in_n313) );
  OAI2BB2X1 reg_in_U575 ( .B0(reg_in_n235), .B1(reg_in_n879), .A0N(Din[52]), 
        .A1N(reg_in_n250), .Y(reg_in_n312) );
  OAI2BB2X1 reg_in_U574 ( .B0(reg_in_n235), .B1(reg_in_n911), .A0N(Din[51]), 
        .A1N(reg_in_n251), .Y(reg_in_n311) );
  OAI2BB2X1 reg_in_U573 ( .B0(reg_in_n235), .B1(reg_in_n943), .A0N(Din[50]), 
        .A1N(reg_in_n251), .Y(reg_in_n310) );
  OAI2BB2X1 reg_in_U572 ( .B0(reg_in_n235), .B1(reg_in_n975), .A0N(Din[49]), 
        .A1N(reg_in_n251), .Y(reg_in_n309) );
  OAI2BB2X1 reg_in_U571 ( .B0(reg_in_n234), .B1(reg_in_n1007), .A0N(Din[48]), 
        .A1N(reg_in_n251), .Y(reg_in_n308) );
  OAI2BB2X1 reg_in_U570 ( .B0(reg_in_n234), .B1(reg_in_n782), .A0N(Din[47]), 
        .A1N(reg_in_n251), .Y(reg_in_n307) );
  OAI2BB2X1 reg_in_U569 ( .B0(reg_in_n234), .B1(reg_in_n814), .A0N(Din[46]), 
        .A1N(reg_in_n251), .Y(reg_in_n306) );
  OAI2BB2X1 reg_in_U568 ( .B0(reg_in_n234), .B1(reg_in_n846), .A0N(Din[45]), 
        .A1N(reg_in_n252), .Y(reg_in_n305) );
  OAI2BB2X1 reg_in_U567 ( .B0(reg_in_n234), .B1(reg_in_n878), .A0N(Din[44]), 
        .A1N(reg_in_n252), .Y(reg_in_n304) );
  OAI2BB2X1 reg_in_U566 ( .B0(reg_in_n234), .B1(reg_in_n910), .A0N(Din[43]), 
        .A1N(reg_in_n252), .Y(reg_in_n303) );
  OAI2BB2X1 reg_in_U565 ( .B0(reg_in_n234), .B1(reg_in_n942), .A0N(Din[42]), 
        .A1N(reg_in_n252), .Y(reg_in_n302) );
  OAI2BB2X1 reg_in_U564 ( .B0(reg_in_n249), .B1(reg_in_n974), .A0N(Din[41]), 
        .A1N(reg_in_n252), .Y(reg_in_n301) );
  OAI2BB2X1 reg_in_U563 ( .B0(reg_in_n248), .B1(reg_in_n1006), .A0N(Din[40]), 
        .A1N(reg_in_n252), .Y(reg_in_n300) );
  OAI2BB2X1 reg_in_U562 ( .B0(reg_in_n241), .B1(reg_in_n781), .A0N(Din[39]), 
        .A1N(reg_in_n253), .Y(reg_in_n299) );
  OAI2BB2X1 reg_in_U561 ( .B0(reg_in_n251), .B1(reg_in_n813), .A0N(Din[38]), 
        .A1N(reg_in_n253), .Y(reg_in_n298) );
  OAI2BB2X1 reg_in_U560 ( .B0(reg_in_n250), .B1(reg_in_n845), .A0N(Din[37]), 
        .A1N(reg_in_n253), .Y(reg_in_n297) );
  OAI2BB2X1 reg_in_U559 ( .B0(reg_in_n235), .B1(reg_in_n877), .A0N(Din[36]), 
        .A1N(reg_in_n252), .Y(reg_in_n296) );
  OAI2BB2X1 reg_in_U558 ( .B0(reg_in_n240), .B1(reg_in_n909), .A0N(Din[35]), 
        .A1N(reg_in_n252), .Y(reg_in_n295) );
  OAI2BB2X1 reg_in_U557 ( .B0(reg_in_n249), .B1(reg_in_n941), .A0N(Din[34]), 
        .A1N(reg_in_n240), .Y(reg_in_n294) );
  OAI2BB2X1 reg_in_U556 ( .B0(reg_in_n248), .B1(reg_in_n973), .A0N(Din[33]), 
        .A1N(reg_in_n252), .Y(reg_in_n293) );
  OAI2BB2X1 reg_in_U555 ( .B0(reg_in_n241), .B1(reg_in_n1005), .A0N(Din[32]), 
        .A1N(reg_in_n240), .Y(reg_in_n292) );
  OAI2BB2X1 reg_in_U554 ( .B0(reg_in_n234), .B1(reg_in_n780), .A0N(Din[31]), 
        .A1N(reg_in_n240), .Y(reg_in_n291) );
  OAI2BB2X1 reg_in_U553 ( .B0(reg_in_n234), .B1(reg_in_n812), .A0N(Din[30]), 
        .A1N(reg_in_n240), .Y(reg_in_n290) );
  OAI2BB2X1 reg_in_U552 ( .B0(reg_in_n234), .B1(reg_in_n844), .A0N(Din[29]), 
        .A1N(reg_in_n240), .Y(reg_in_n289) );
  OAI2BB2X1 reg_in_U551 ( .B0(reg_in_n234), .B1(reg_in_n876), .A0N(Din[28]), 
        .A1N(reg_in_n241), .Y(reg_in_n288) );
  OAI2BB2X1 reg_in_U550 ( .B0(reg_in_n234), .B1(reg_in_n908), .A0N(Din[27]), 
        .A1N(reg_in_n241), .Y(reg_in_n287) );
  OAI2BB2X1 reg_in_U549 ( .B0(reg_in_n235), .B1(reg_in_n940), .A0N(Din[26]), 
        .A1N(reg_in_n241), .Y(reg_in_n286) );
  OAI2BB2X1 reg_in_U548 ( .B0(reg_in_n235), .B1(reg_in_n972), .A0N(Din[25]), 
        .A1N(reg_in_n242), .Y(reg_in_n285) );
  OAI2BB2X1 reg_in_U547 ( .B0(reg_in_n235), .B1(reg_in_n1004), .A0N(Din[24]), 
        .A1N(reg_in_n242), .Y(reg_in_n284) );
  OAI2BB2X1 reg_in_U546 ( .B0(reg_in_n235), .B1(reg_in_n779), .A0N(Din[23]), 
        .A1N(reg_in_n242), .Y(reg_in_n283) );
  OAI2BB2X1 reg_in_U545 ( .B0(reg_in_n238), .B1(reg_in_n811), .A0N(Din[22]), 
        .A1N(reg_in_n242), .Y(reg_in_n282) );
  OAI2BB2X1 reg_in_U544 ( .B0(reg_in_n236), .B1(reg_in_n843), .A0N(Din[21]), 
        .A1N(reg_in_n243), .Y(reg_in_n281) );
  OAI2BB2X1 reg_in_U543 ( .B0(reg_in_n236), .B1(reg_in_n875), .A0N(Din[20]), 
        .A1N(reg_in_n243), .Y(reg_in_n280) );
  OAI2BB2X1 reg_in_U542 ( .B0(reg_in_n236), .B1(reg_in_n907), .A0N(Din[19]), 
        .A1N(reg_in_n243), .Y(reg_in_n279) );
  OAI2BB2X1 reg_in_U541 ( .B0(reg_in_n236), .B1(reg_in_n939), .A0N(Din[18]), 
        .A1N(reg_in_n243), .Y(reg_in_n278) );
  OAI2BB2X1 reg_in_U540 ( .B0(reg_in_n236), .B1(reg_in_n971), .A0N(Din[17]), 
        .A1N(reg_in_n244), .Y(reg_in_n277) );
  OAI2BB2X1 reg_in_U539 ( .B0(reg_in_n237), .B1(reg_in_n1003), .A0N(Din[16]), 
        .A1N(reg_in_n244), .Y(reg_in_n276) );
  OAI2BB2X1 reg_in_U538 ( .B0(reg_in_n237), .B1(reg_in_n778), .A0N(Din[15]), 
        .A1N(reg_in_n244), .Y(reg_in_n275) );
  OAI2BB2X1 reg_in_U537 ( .B0(reg_in_n237), .B1(reg_in_n810), .A0N(Din[14]), 
        .A1N(reg_in_n244), .Y(reg_in_n274) );
  OAI2BB2X1 reg_in_U536 ( .B0(reg_in_n237), .B1(reg_in_n842), .A0N(Din[13]), 
        .A1N(reg_in_n245), .Y(reg_in_n273) );
  OAI2BB2X1 reg_in_U535 ( .B0(reg_in_n237), .B1(reg_in_n874), .A0N(Din[12]), 
        .A1N(reg_in_n245), .Y(reg_in_n272) );
  OAI2BB2X1 reg_in_U534 ( .B0(reg_in_n238), .B1(reg_in_n906), .A0N(Din[11]), 
        .A1N(reg_in_n252), .Y(reg_in_n271) );
  OAI2BB2X1 reg_in_U533 ( .B0(reg_in_n238), .B1(reg_in_n938), .A0N(Din[10]), 
        .A1N(reg_in_n244), .Y(reg_in_n270) );
  OAI2BB2X1 reg_in_U532 ( .B0(reg_in_n238), .B1(reg_in_n970), .A0N(Din[9]), 
        .A1N(reg_in_n244), .Y(reg_in_n269) );
  OAI2BB2X1 reg_in_U531 ( .B0(reg_in_n239), .B1(reg_in_n1002), .A0N(Din[8]), 
        .A1N(reg_in_n243), .Y(reg_in_n268) );
  OAI2BB2X1 reg_in_U530 ( .B0(reg_in_n247), .B1(reg_in_n777), .A0N(Din[7]), 
        .A1N(reg_in_n243), .Y(reg_in_n267) );
  OAI2BB2X1 reg_in_U529 ( .B0(reg_in_n246), .B1(reg_in_n809), .A0N(Din[6]), 
        .A1N(reg_in_n242), .Y(reg_in_n266) );
  OAI2BB2X1 reg_in_U528 ( .B0(reg_in_n243), .B1(reg_in_n841), .A0N(Din[5]), 
        .A1N(reg_in_n242), .Y(reg_in_n265) );
  OAI2BB2X1 reg_in_U527 ( .B0(reg_in_n239), .B1(reg_in_n873), .A0N(Din[4]), 
        .A1N(reg_in_n241), .Y(reg_in_n264) );
  OAI2BB2X1 reg_in_U526 ( .B0(reg_in_n239), .B1(reg_in_n905), .A0N(Din[3]), 
        .A1N(reg_in_n241), .Y(reg_in_n263) );
  OAI2BB2X1 reg_in_U525 ( .B0(reg_in_n238), .B1(reg_in_n937), .A0N(Din[2]), 
        .A1N(reg_in_n240), .Y(reg_in_n262) );
  OAI2BB2X1 reg_in_U524 ( .B0(reg_in_n239), .B1(reg_in_n969), .A0N(Din[1]), 
        .A1N(reg_in_n252), .Y(reg_in_n261) );
  OAI2BB2X1 reg_in_U523 ( .B0(reg_in_n238), .B1(reg_in_n1001), .A0N(Din[0]), 
        .A1N(reg_in_n245), .Y(reg_in_n260) );
  NAND2BX1 reg_in_U522 ( .AN(reg_in_pf0), .B(reg_in_pf1), .Y(reg_in_n1) );
  NAND2BX1 reg_in_U521 ( .AN(reg_in_pbv0), .B(reg_in_pbv1), .Y(reg_in_n258) );
  OAI2BB2X1 reg_in_U520 ( .B0(reg_in_n2), .B1(reg_in_n777), .A0N(
        plain_byte_in[7]), .A1N(reg_in_n21), .Y(reg_in_n771) );
  OAI2BB2X1 reg_in_U519 ( .B0(reg_in_n2), .B1(reg_in_n809), .A0N(
        plain_byte_in[6]), .A1N(reg_in_n180), .Y(reg_in_n739) );
  OAI2BB2X1 reg_in_U518 ( .B0(reg_in_n2), .B1(reg_in_n841), .A0N(
        plain_byte_in[5]), .A1N(reg_in_n21), .Y(reg_in_n707) );
  OAI2BB2X1 reg_in_U517 ( .B0(reg_in_n2), .B1(reg_in_n873), .A0N(
        plain_byte_in[4]), .A1N(reg_in_n21), .Y(reg_in_n675) );
  OAI2BB2X1 reg_in_U516 ( .B0(reg_in_n2), .B1(reg_in_n905), .A0N(
        plain_byte_in[3]), .A1N(reg_in_n179), .Y(reg_in_n643) );
  OAI2BB2X1 reg_in_U515 ( .B0(reg_in_n2), .B1(reg_in_n937), .A0N(
        plain_byte_in[2]), .A1N(reg_in_n21), .Y(reg_in_n611) );
  OAI2BB2X1 reg_in_U514 ( .B0(reg_in_n2), .B1(reg_in_n969), .A0N(
        plain_byte_in[1]), .A1N(reg_in_n21), .Y(reg_in_n579) );
  OAI2BB2X1 reg_in_U513 ( .B0(reg_in_n2), .B1(reg_in_n1001), .A0N(
        plain_byte_in[0]), .A1N(reg_in_n171), .Y(reg_in_n547) );
  INVX1 reg_in_U512 ( .A(reg_in_n1), .Y(reg_in_n219) );
  INVX1 reg_in_U511 ( .A(reg_in_n258), .Y(reg_in_n216) );
  INVX1 reg_in_U510 ( .A(reg_in_n258), .Y(reg_in_n215) );
  INVX1 reg_in_U509 ( .A(reg_in_n258), .Y(reg_in_n214) );
  INVX1 reg_in_U508 ( .A(reg_in_n258), .Y(reg_in_n213) );
  INVX1 reg_in_U507 ( .A(reg_in_n258), .Y(reg_in_n212) );
  INVX1 reg_in_U506 ( .A(reg_in_n258), .Y(reg_in_n211) );
  INVX1 reg_in_U505 ( .A(reg_in_n258), .Y(reg_in_n210) );
  OAI22X1 reg_in_U504 ( .A0(reg_in_n807), .A1(reg_in_n37), .B0(reg_in_n12), 
        .B1(reg_in_n808), .Y(reg_in_n740) );
  OAI22X1 reg_in_U503 ( .A0(reg_in_n839), .A1(reg_in_n50), .B0(reg_in_n12), 
        .B1(reg_in_n840), .Y(reg_in_n708) );
  OAI22X1 reg_in_U502 ( .A0(reg_in_n871), .A1(reg_in_n65), .B0(reg_in_n15), 
        .B1(reg_in_n872), .Y(reg_in_n676) );
  OAI22X1 reg_in_U501 ( .A0(reg_in_n903), .A1(reg_in_n79), .B0(reg_in_n3), 
        .B1(reg_in_n904), .Y(reg_in_n644) );
  OAI22X1 reg_in_U500 ( .A0(reg_in_n935), .A1(reg_in_n93), .B0(reg_in_n10), 
        .B1(reg_in_n936), .Y(reg_in_n612) );
  OAI22X1 reg_in_U499 ( .A0(reg_in_n967), .A1(reg_in_n107), .B0(reg_in_n7), 
        .B1(reg_in_n968), .Y(reg_in_n580) );
  OAI22X1 reg_in_U498 ( .A0(reg_in_n999), .A1(reg_in_n124), .B0(reg_in_n5), 
        .B1(reg_in_n1000), .Y(reg_in_n548) );
  OAI22X1 reg_in_U497 ( .A0(reg_in_n1031), .A1(reg_in_n116), .B0(reg_in_n7), 
        .B1(reg_in_n1032), .Y(reg_in_n516) );
  OAI22X1 reg_in_U496 ( .A0(reg_in_n777), .A1(reg_in_n22), .B0(reg_in_n21), 
        .B1(reg_in_n778), .Y(reg_in_n770) );
  OAI22X1 reg_in_U495 ( .A0(reg_in_n778), .A1(reg_in_n22), .B0(reg_in_n7), 
        .B1(reg_in_n779), .Y(reg_in_n769) );
  OAI22X1 reg_in_U494 ( .A0(reg_in_n779), .A1(reg_in_n23), .B0(reg_in_n20), 
        .B1(reg_in_n780), .Y(reg_in_n768) );
  OAI22X1 reg_in_U493 ( .A0(reg_in_n780), .A1(reg_in_n23), .B0(reg_in_n21), 
        .B1(reg_in_n781), .Y(reg_in_n767) );
  OAI22X1 reg_in_U492 ( .A0(reg_in_n781), .A1(reg_in_n24), .B0(reg_in_n21), 
        .B1(reg_in_n782), .Y(reg_in_n766) );
  OAI22X1 reg_in_U491 ( .A0(reg_in_n782), .A1(reg_in_n24), .B0(reg_in_n2), 
        .B1(reg_in_n783), .Y(reg_in_n765) );
  OAI22X1 reg_in_U490 ( .A0(reg_in_n783), .A1(reg_in_n25), .B0(reg_in_n17), 
        .B1(reg_in_n784), .Y(reg_in_n764) );
  OAI22X1 reg_in_U489 ( .A0(reg_in_n784), .A1(reg_in_n25), .B0(reg_in_n20), 
        .B1(reg_in_n785), .Y(reg_in_n763) );
  OAI22X1 reg_in_U488 ( .A0(reg_in_n785), .A1(reg_in_n26), .B0(reg_in_n21), 
        .B1(reg_in_n786), .Y(reg_in_n762) );
  OAI22X1 reg_in_U487 ( .A0(reg_in_n786), .A1(reg_in_n26), .B0(reg_in_n21), 
        .B1(reg_in_n787), .Y(reg_in_n761) );
  OAI22X1 reg_in_U486 ( .A0(reg_in_n787), .A1(reg_in_n27), .B0(reg_in_n21), 
        .B1(reg_in_n788), .Y(reg_in_n760) );
  OAI22X1 reg_in_U485 ( .A0(reg_in_n788), .A1(reg_in_n27), .B0(reg_in_n21), 
        .B1(reg_in_n789), .Y(reg_in_n759) );
  OAI22X1 reg_in_U484 ( .A0(reg_in_n789), .A1(reg_in_n28), .B0(reg_in_n21), 
        .B1(reg_in_n790), .Y(reg_in_n758) );
  OAI22X1 reg_in_U483 ( .A0(reg_in_n790), .A1(reg_in_n28), .B0(reg_in_n3), 
        .B1(reg_in_n791), .Y(reg_in_n757) );
  OAI22X1 reg_in_U482 ( .A0(reg_in_n791), .A1(reg_in_n29), .B0(reg_in_n12), 
        .B1(reg_in_n792), .Y(reg_in_n756) );
  OAI22X1 reg_in_U481 ( .A0(reg_in_n792), .A1(reg_in_n29), .B0(reg_in_n17), 
        .B1(reg_in_n793), .Y(reg_in_n755) );
  OAI22X1 reg_in_U480 ( .A0(reg_in_n793), .A1(reg_in_n30), .B0(reg_in_n19), 
        .B1(reg_in_n794), .Y(reg_in_n754) );
  OAI22X1 reg_in_U479 ( .A0(reg_in_n794), .A1(reg_in_n30), .B0(reg_in_n20), 
        .B1(reg_in_n795), .Y(reg_in_n753) );
  OAI22X1 reg_in_U478 ( .A0(reg_in_n795), .A1(reg_in_n31), .B0(reg_in_n20), 
        .B1(reg_in_n796), .Y(reg_in_n752) );
  OAI22X1 reg_in_U477 ( .A0(reg_in_n796), .A1(reg_in_n31), .B0(reg_in_n21), 
        .B1(reg_in_n797), .Y(reg_in_n751) );
  OAI22X1 reg_in_U476 ( .A0(reg_in_n797), .A1(reg_in_n32), .B0(reg_in_n20), 
        .B1(reg_in_n798), .Y(reg_in_n750) );
  OAI22X1 reg_in_U475 ( .A0(reg_in_n798), .A1(reg_in_n32), .B0(reg_in_n20), 
        .B1(reg_in_n799), .Y(reg_in_n749) );
  OAI22X1 reg_in_U474 ( .A0(reg_in_n799), .A1(reg_in_n33), .B0(reg_in_n20), 
        .B1(reg_in_n800), .Y(reg_in_n748) );
  OAI22X1 reg_in_U473 ( .A0(reg_in_n800), .A1(reg_in_n33), .B0(reg_in_n20), 
        .B1(reg_in_n801), .Y(reg_in_n747) );
  OAI22X1 reg_in_U472 ( .A0(reg_in_n801), .A1(reg_in_n34), .B0(reg_in_n20), 
        .B1(reg_in_n802), .Y(reg_in_n746) );
  OAI22X1 reg_in_U471 ( .A0(reg_in_n802), .A1(reg_in_n34), .B0(reg_in_n20), 
        .B1(reg_in_n803), .Y(reg_in_n745) );
  OAI22X1 reg_in_U470 ( .A0(reg_in_n803), .A1(reg_in_n35), .B0(reg_in_n20), 
        .B1(reg_in_n804), .Y(reg_in_n744) );
  OAI22X1 reg_in_U469 ( .A0(reg_in_n804), .A1(reg_in_n35), .B0(reg_in_n20), 
        .B1(reg_in_n805), .Y(reg_in_n743) );
  OAI22X1 reg_in_U468 ( .A0(reg_in_n805), .A1(reg_in_n36), .B0(reg_in_n20), 
        .B1(reg_in_n806), .Y(reg_in_n742) );
  OAI22X1 reg_in_U467 ( .A0(reg_in_n806), .A1(reg_in_n36), .B0(reg_in_n3), 
        .B1(reg_in_n807), .Y(reg_in_n741) );
  OAI22X1 reg_in_U466 ( .A0(reg_in_n809), .A1(reg_in_n38), .B0(reg_in_n17), 
        .B1(reg_in_n810), .Y(reg_in_n738) );
  OAI22X1 reg_in_U465 ( .A0(reg_in_n810), .A1(reg_in_n37), .B0(reg_in_n17), 
        .B1(reg_in_n811), .Y(reg_in_n737) );
  OAI22X1 reg_in_U464 ( .A0(reg_in_n811), .A1(reg_in_n37), .B0(reg_in_n19), 
        .B1(reg_in_n812), .Y(reg_in_n736) );
  OAI22X1 reg_in_U463 ( .A0(reg_in_n812), .A1(reg_in_n38), .B0(reg_in_n19), 
        .B1(reg_in_n813), .Y(reg_in_n735) );
  OAI22X1 reg_in_U462 ( .A0(reg_in_n813), .A1(reg_in_n38), .B0(reg_in_n19), 
        .B1(reg_in_n814), .Y(reg_in_n734) );
  OAI22X1 reg_in_U461 ( .A0(reg_in_n814), .A1(reg_in_n39), .B0(reg_in_n19), 
        .B1(reg_in_n815), .Y(reg_in_n733) );
  OAI22X1 reg_in_U460 ( .A0(reg_in_n815), .A1(reg_in_n40), .B0(reg_in_n19), 
        .B1(reg_in_n816), .Y(reg_in_n732) );
  OAI22X1 reg_in_U459 ( .A0(reg_in_n816), .A1(reg_in_n39), .B0(reg_in_n19), 
        .B1(reg_in_n817), .Y(reg_in_n731) );
  OAI22X1 reg_in_U458 ( .A0(reg_in_n817), .A1(reg_in_n39), .B0(reg_in_n19), 
        .B1(reg_in_n818), .Y(reg_in_n730) );
  OAI22X1 reg_in_U457 ( .A0(reg_in_n818), .A1(reg_in_n40), .B0(reg_in_n19), 
        .B1(reg_in_n819), .Y(reg_in_n729) );
  OAI22X1 reg_in_U456 ( .A0(reg_in_n819), .A1(reg_in_n40), .B0(reg_in_n19), 
        .B1(reg_in_n820), .Y(reg_in_n728) );
  OAI22X1 reg_in_U455 ( .A0(reg_in_n820), .A1(reg_in_n41), .B0(reg_in_n19), 
        .B1(reg_in_n821), .Y(reg_in_n727) );
  OAI22X1 reg_in_U454 ( .A0(reg_in_n821), .A1(reg_in_n41), .B0(reg_in_n19), 
        .B1(reg_in_n822), .Y(reg_in_n726) );
  OAI22X1 reg_in_U453 ( .A0(reg_in_n822), .A1(reg_in_n42), .B0(reg_in_n19), 
        .B1(reg_in_n823), .Y(reg_in_n725) );
  OAI22X1 reg_in_U452 ( .A0(reg_in_n823), .A1(reg_in_n42), .B0(reg_in_n18), 
        .B1(reg_in_n824), .Y(reg_in_n724) );
  OAI22X1 reg_in_U451 ( .A0(reg_in_n824), .A1(reg_in_n43), .B0(reg_in_n18), 
        .B1(reg_in_n825), .Y(reg_in_n723) );
  OAI22X1 reg_in_U450 ( .A0(reg_in_n825), .A1(reg_in_n43), .B0(reg_in_n18), 
        .B1(reg_in_n826), .Y(reg_in_n722) );
  OAI22X1 reg_in_U449 ( .A0(reg_in_n826), .A1(reg_in_n44), .B0(reg_in_n18), 
        .B1(reg_in_n827), .Y(reg_in_n721) );
  OAI22X1 reg_in_U448 ( .A0(reg_in_n827), .A1(reg_in_n44), .B0(reg_in_n18), 
        .B1(reg_in_n828), .Y(reg_in_n720) );
  OAI22X1 reg_in_U447 ( .A0(reg_in_n828), .A1(reg_in_n45), .B0(reg_in_n18), 
        .B1(reg_in_n829), .Y(reg_in_n719) );
  OAI22X1 reg_in_U446 ( .A0(reg_in_n829), .A1(reg_in_n45), .B0(reg_in_n18), 
        .B1(reg_in_n830), .Y(reg_in_n718) );
  OAI22X1 reg_in_U445 ( .A0(reg_in_n830), .A1(reg_in_n46), .B0(reg_in_n18), 
        .B1(reg_in_n831), .Y(reg_in_n717) );
  OAI22X1 reg_in_U444 ( .A0(reg_in_n831), .A1(reg_in_n46), .B0(reg_in_n18), 
        .B1(reg_in_n832), .Y(reg_in_n716) );
  OAI22X1 reg_in_U443 ( .A0(reg_in_n832), .A1(reg_in_n47), .B0(reg_in_n18), 
        .B1(reg_in_n833), .Y(reg_in_n715) );
  OAI22X1 reg_in_U442 ( .A0(reg_in_n833), .A1(reg_in_n47), .B0(reg_in_n18), 
        .B1(reg_in_n834), .Y(reg_in_n714) );
  OAI22X1 reg_in_U441 ( .A0(reg_in_n834), .A1(reg_in_n48), .B0(reg_in_n18), 
        .B1(reg_in_n835), .Y(reg_in_n713) );
  OAI22X1 reg_in_U440 ( .A0(reg_in_n835), .A1(reg_in_n48), .B0(reg_in_n18), 
        .B1(reg_in_n836), .Y(reg_in_n712) );
  OAI22X1 reg_in_U439 ( .A0(reg_in_n836), .A1(reg_in_n49), .B0(reg_in_n17), 
        .B1(reg_in_n837), .Y(reg_in_n711) );
  OAI22X1 reg_in_U438 ( .A0(reg_in_n837), .A1(reg_in_n49), .B0(reg_in_n2), 
        .B1(reg_in_n838), .Y(reg_in_n710) );
  OAI22X1 reg_in_U437 ( .A0(reg_in_n838), .A1(reg_in_n50), .B0(reg_in_n2), 
        .B1(reg_in_n839), .Y(reg_in_n709) );
  OAI22X1 reg_in_U436 ( .A0(reg_in_n841), .A1(reg_in_n51), .B0(reg_in_n13), 
        .B1(reg_in_n842), .Y(reg_in_n706) );
  OAI22X1 reg_in_U435 ( .A0(reg_in_n842), .A1(reg_in_n51), .B0(reg_in_n17), 
        .B1(reg_in_n843), .Y(reg_in_n705) );
  OAI22X1 reg_in_U434 ( .A0(reg_in_n843), .A1(reg_in_n52), .B0(reg_in_n17), 
        .B1(reg_in_n844), .Y(reg_in_n704) );
  OAI22X1 reg_in_U433 ( .A0(reg_in_n844), .A1(reg_in_n52), .B0(reg_in_n17), 
        .B1(reg_in_n845), .Y(reg_in_n703) );
  OAI22X1 reg_in_U432 ( .A0(reg_in_n845), .A1(reg_in_n53), .B0(reg_in_n17), 
        .B1(reg_in_n846), .Y(reg_in_n702) );
  OAI22X1 reg_in_U431 ( .A0(reg_in_n846), .A1(reg_in_n53), .B0(reg_in_n17), 
        .B1(reg_in_n847), .Y(reg_in_n701) );
  OAI22X1 reg_in_U430 ( .A0(reg_in_n847), .A1(reg_in_n54), .B0(reg_in_n17), 
        .B1(reg_in_n848), .Y(reg_in_n700) );
  OAI22X1 reg_in_U429 ( .A0(reg_in_n848), .A1(reg_in_n54), .B0(reg_in_n17), 
        .B1(reg_in_n849), .Y(reg_in_n699) );
  OAI22X1 reg_in_U428 ( .A0(reg_in_n849), .A1(reg_in_n55), .B0(reg_in_n16), 
        .B1(reg_in_n850), .Y(reg_in_n698) );
  OAI22X1 reg_in_U427 ( .A0(reg_in_n850), .A1(reg_in_n55), .B0(reg_in_n16), 
        .B1(reg_in_n851), .Y(reg_in_n697) );
  OAI22X1 reg_in_U426 ( .A0(reg_in_n851), .A1(reg_in_n56), .B0(reg_in_n16), 
        .B1(reg_in_n852), .Y(reg_in_n696) );
  OAI22X1 reg_in_U425 ( .A0(reg_in_n852), .A1(reg_in_n56), .B0(reg_in_n16), 
        .B1(reg_in_n853), .Y(reg_in_n695) );
  OAI22X1 reg_in_U424 ( .A0(reg_in_n853), .A1(reg_in_n57), .B0(reg_in_n16), 
        .B1(reg_in_n854), .Y(reg_in_n694) );
  OAI22X1 reg_in_U423 ( .A0(reg_in_n854), .A1(reg_in_n57), .B0(reg_in_n16), 
        .B1(reg_in_n855), .Y(reg_in_n693) );
  OAI22X1 reg_in_U422 ( .A0(reg_in_n855), .A1(reg_in_n58), .B0(reg_in_n16), 
        .B1(reg_in_n856), .Y(reg_in_n692) );
  OAI22X1 reg_in_U421 ( .A0(reg_in_n856), .A1(reg_in_n58), .B0(reg_in_n16), 
        .B1(reg_in_n857), .Y(reg_in_n691) );
  OAI22X1 reg_in_U420 ( .A0(reg_in_n857), .A1(reg_in_n59), .B0(reg_in_n16), 
        .B1(reg_in_n858), .Y(reg_in_n690) );
  OAI22X1 reg_in_U419 ( .A0(reg_in_n858), .A1(reg_in_n59), .B0(reg_in_n16), 
        .B1(reg_in_n859), .Y(reg_in_n689) );
  OAI22X1 reg_in_U418 ( .A0(reg_in_n859), .A1(reg_in_n60), .B0(reg_in_n16), 
        .B1(reg_in_n860), .Y(reg_in_n688) );
  OAI22X1 reg_in_U417 ( .A0(reg_in_n860), .A1(reg_in_n60), .B0(reg_in_n16), 
        .B1(reg_in_n861), .Y(reg_in_n687) );
  OAI22X1 reg_in_U416 ( .A0(reg_in_n861), .A1(reg_in_n61), .B0(reg_in_n16), 
        .B1(reg_in_n862), .Y(reg_in_n686) );
  OAI22X1 reg_in_U415 ( .A0(reg_in_n862), .A1(reg_in_n61), .B0(reg_in_n15), 
        .B1(reg_in_n863), .Y(reg_in_n685) );
  OAI22X1 reg_in_U414 ( .A0(reg_in_n863), .A1(reg_in_n62), .B0(reg_in_n15), 
        .B1(reg_in_n864), .Y(reg_in_n684) );
  OAI22X1 reg_in_U413 ( .A0(reg_in_n864), .A1(reg_in_n62), .B0(reg_in_n15), 
        .B1(reg_in_n865), .Y(reg_in_n683) );
  OAI22X1 reg_in_U412 ( .A0(reg_in_n865), .A1(reg_in_n63), .B0(reg_in_n15), 
        .B1(reg_in_n866), .Y(reg_in_n682) );
  OAI22X1 reg_in_U411 ( .A0(reg_in_n866), .A1(reg_in_n63), .B0(reg_in_n15), 
        .B1(reg_in_n867), .Y(reg_in_n681) );
  OAI22X1 reg_in_U410 ( .A0(reg_in_n867), .A1(reg_in_n64), .B0(reg_in_n15), 
        .B1(reg_in_n868), .Y(reg_in_n680) );
  OAI22X1 reg_in_U409 ( .A0(reg_in_n868), .A1(reg_in_n64), .B0(reg_in_n15), 
        .B1(reg_in_n869), .Y(reg_in_n679) );
  OAI22X1 reg_in_U408 ( .A0(reg_in_n869), .A1(reg_in_n65), .B0(reg_in_n15), 
        .B1(reg_in_n870), .Y(reg_in_n678) );
  OAI22X1 reg_in_U407 ( .A0(reg_in_n870), .A1(reg_in_n65), .B0(reg_in_n15), 
        .B1(reg_in_n871), .Y(reg_in_n677) );
  OAI22X1 reg_in_U406 ( .A0(reg_in_n873), .A1(reg_in_n66), .B0(reg_in_n15), 
        .B1(reg_in_n874), .Y(reg_in_n674) );
  OAI22X1 reg_in_U405 ( .A0(reg_in_n874), .A1(reg_in_n66), .B0(reg_in_n14), 
        .B1(reg_in_n875), .Y(reg_in_n673) );
  OAI22X1 reg_in_U404 ( .A0(reg_in_n875), .A1(reg_in_n66), .B0(reg_in_n14), 
        .B1(reg_in_n876), .Y(reg_in_n672) );
  OAI22X1 reg_in_U403 ( .A0(reg_in_n876), .A1(reg_in_n67), .B0(reg_in_n14), 
        .B1(reg_in_n877), .Y(reg_in_n671) );
  OAI22X1 reg_in_U402 ( .A0(reg_in_n877), .A1(reg_in_n67), .B0(reg_in_n14), 
        .B1(reg_in_n878), .Y(reg_in_n670) );
  OAI22X1 reg_in_U401 ( .A0(reg_in_n878), .A1(reg_in_n68), .B0(reg_in_n14), 
        .B1(reg_in_n879), .Y(reg_in_n669) );
  OAI22X1 reg_in_U400 ( .A0(reg_in_n879), .A1(reg_in_n68), .B0(reg_in_n14), 
        .B1(reg_in_n880), .Y(reg_in_n668) );
  OAI22X1 reg_in_U399 ( .A0(reg_in_n880), .A1(reg_in_n69), .B0(reg_in_n14), 
        .B1(reg_in_n881), .Y(reg_in_n667) );
  OAI22X1 reg_in_U398 ( .A0(reg_in_n881), .A1(reg_in_n69), .B0(reg_in_n14), 
        .B1(reg_in_n882), .Y(reg_in_n666) );
  OAI22X1 reg_in_U397 ( .A0(reg_in_n882), .A1(reg_in_n70), .B0(reg_in_n14), 
        .B1(reg_in_n883), .Y(reg_in_n665) );
  OAI22X1 reg_in_U396 ( .A0(reg_in_n883), .A1(reg_in_n70), .B0(reg_in_n14), 
        .B1(reg_in_n884), .Y(reg_in_n664) );
  OAI22X1 reg_in_U395 ( .A0(reg_in_n884), .A1(reg_in_n71), .B0(reg_in_n14), 
        .B1(reg_in_n885), .Y(reg_in_n663) );
  OAI22X1 reg_in_U394 ( .A0(reg_in_n885), .A1(reg_in_n71), .B0(reg_in_n14), 
        .B1(reg_in_n886), .Y(reg_in_n662) );
  OAI22X1 reg_in_U393 ( .A0(reg_in_n886), .A1(reg_in_n72), .B0(reg_in_n14), 
        .B1(reg_in_n887), .Y(reg_in_n661) );
  OAI22X1 reg_in_U392 ( .A0(reg_in_n887), .A1(reg_in_n72), .B0(reg_in_n13), 
        .B1(reg_in_n888), .Y(reg_in_n660) );
  OAI22X1 reg_in_U391 ( .A0(reg_in_n888), .A1(reg_in_n73), .B0(reg_in_n13), 
        .B1(reg_in_n889), .Y(reg_in_n659) );
  OAI22X1 reg_in_U390 ( .A0(reg_in_n889), .A1(reg_in_n73), .B0(reg_in_n13), 
        .B1(reg_in_n890), .Y(reg_in_n658) );
  OAI22X1 reg_in_U389 ( .A0(reg_in_n890), .A1(reg_in_n74), .B0(reg_in_n13), 
        .B1(reg_in_n891), .Y(reg_in_n657) );
  OAI22X1 reg_in_U388 ( .A0(reg_in_n891), .A1(reg_in_n74), .B0(reg_in_n13), 
        .B1(reg_in_n892), .Y(reg_in_n656) );
  OAI22X1 reg_in_U387 ( .A0(reg_in_n892), .A1(reg_in_n75), .B0(reg_in_n13), 
        .B1(reg_in_n893), .Y(reg_in_n655) );
  OAI22X1 reg_in_U386 ( .A0(reg_in_n893), .A1(reg_in_n75), .B0(reg_in_n13), 
        .B1(reg_in_n894), .Y(reg_in_n654) );
  OAI22X1 reg_in_U385 ( .A0(reg_in_n894), .A1(reg_in_n76), .B0(reg_in_n13), 
        .B1(reg_in_n895), .Y(reg_in_n653) );
  OAI22X1 reg_in_U384 ( .A0(reg_in_n895), .A1(reg_in_n76), .B0(reg_in_n13), 
        .B1(reg_in_n896), .Y(reg_in_n652) );
  OAI22X1 reg_in_U383 ( .A0(reg_in_n896), .A1(reg_in_n77), .B0(reg_in_n13), 
        .B1(reg_in_n897), .Y(reg_in_n651) );
  OAI22X1 reg_in_U382 ( .A0(reg_in_n897), .A1(reg_in_n77), .B0(reg_in_n13), 
        .B1(reg_in_n898), .Y(reg_in_n650) );
  OAI22X1 reg_in_U381 ( .A0(reg_in_n898), .A1(reg_in_n78), .B0(reg_in_n13), 
        .B1(reg_in_n899), .Y(reg_in_n649) );
  OAI22X1 reg_in_U380 ( .A0(reg_in_n899), .A1(reg_in_n78), .B0(reg_in_n2), 
        .B1(reg_in_n900), .Y(reg_in_n648) );
  OAI22X1 reg_in_U379 ( .A0(reg_in_n900), .A1(reg_in_n79), .B0(reg_in_n3), 
        .B1(reg_in_n901), .Y(reg_in_n647) );
  OAI22X1 reg_in_U378 ( .A0(reg_in_n901), .A1(reg_in_n79), .B0(reg_in_n7), 
        .B1(reg_in_n902), .Y(reg_in_n646) );
  OAI22X1 reg_in_U377 ( .A0(reg_in_n902), .A1(reg_in_n80), .B0(reg_in_n12), 
        .B1(reg_in_n903), .Y(reg_in_n645) );
  OAI22X1 reg_in_U376 ( .A0(reg_in_n905), .A1(reg_in_n80), .B0(reg_in_n12), 
        .B1(reg_in_n906), .Y(reg_in_n642) );
  OAI22X1 reg_in_U375 ( .A0(reg_in_n906), .A1(reg_in_n80), .B0(reg_in_n12), 
        .B1(reg_in_n907), .Y(reg_in_n641) );
  OAI22X1 reg_in_U374 ( .A0(reg_in_n907), .A1(reg_in_n81), .B0(reg_in_n12), 
        .B1(reg_in_n908), .Y(reg_in_n640) );
  OAI22X1 reg_in_U373 ( .A0(reg_in_n908), .A1(reg_in_n81), .B0(reg_in_n12), 
        .B1(reg_in_n909), .Y(reg_in_n639) );
  OAI22X1 reg_in_U372 ( .A0(reg_in_n909), .A1(reg_in_n82), .B0(reg_in_n12), 
        .B1(reg_in_n910), .Y(reg_in_n638) );
  OAI22X1 reg_in_U371 ( .A0(reg_in_n910), .A1(reg_in_n82), .B0(reg_in_n17), 
        .B1(reg_in_n911), .Y(reg_in_n637) );
  OAI22X1 reg_in_U370 ( .A0(reg_in_n911), .A1(reg_in_n83), .B0(reg_in_n12), 
        .B1(reg_in_n912), .Y(reg_in_n636) );
  OAI22X1 reg_in_U369 ( .A0(reg_in_n912), .A1(reg_in_n83), .B0(reg_in_n11), 
        .B1(reg_in_n913), .Y(reg_in_n635) );
  OAI22X1 reg_in_U368 ( .A0(reg_in_n913), .A1(reg_in_n84), .B0(reg_in_n11), 
        .B1(reg_in_n914), .Y(reg_in_n634) );
  OAI22X1 reg_in_U367 ( .A0(reg_in_n914), .A1(reg_in_n84), .B0(reg_in_n11), 
        .B1(reg_in_n915), .Y(reg_in_n633) );
  OAI22X1 reg_in_U366 ( .A0(reg_in_n915), .A1(reg_in_n85), .B0(reg_in_n11), 
        .B1(reg_in_n916), .Y(reg_in_n632) );
  OAI22X1 reg_in_U365 ( .A0(reg_in_n916), .A1(reg_in_n85), .B0(reg_in_n11), 
        .B1(reg_in_n917), .Y(reg_in_n631) );
  OAI22X1 reg_in_U364 ( .A0(reg_in_n917), .A1(reg_in_n86), .B0(reg_in_n11), 
        .B1(reg_in_n918), .Y(reg_in_n630) );
  OAI22X1 reg_in_U363 ( .A0(reg_in_n918), .A1(reg_in_n86), .B0(reg_in_n11), 
        .B1(reg_in_n919), .Y(reg_in_n629) );
  OAI22X1 reg_in_U362 ( .A0(reg_in_n919), .A1(reg_in_n87), .B0(reg_in_n11), 
        .B1(reg_in_n920), .Y(reg_in_n628) );
  OAI22X1 reg_in_U361 ( .A0(reg_in_n920), .A1(reg_in_n87), .B0(reg_in_n11), 
        .B1(reg_in_n921), .Y(reg_in_n627) );
  OAI22X1 reg_in_U360 ( .A0(reg_in_n921), .A1(reg_in_n88), .B0(reg_in_n11), 
        .B1(reg_in_n922), .Y(reg_in_n626) );
  OAI22X1 reg_in_U359 ( .A0(reg_in_n922), .A1(reg_in_n88), .B0(reg_in_n11), 
        .B1(reg_in_n923), .Y(reg_in_n625) );
  OAI22X1 reg_in_U358 ( .A0(reg_in_n923), .A1(reg_in_n89), .B0(reg_in_n11), 
        .B1(reg_in_n924), .Y(reg_in_n624) );
  OAI22X1 reg_in_U357 ( .A0(reg_in_n924), .A1(reg_in_n89), .B0(reg_in_n11), 
        .B1(reg_in_n925), .Y(reg_in_n623) );
  OAI22X1 reg_in_U356 ( .A0(reg_in_n925), .A1(reg_in_n90), .B0(reg_in_n10), 
        .B1(reg_in_n926), .Y(reg_in_n622) );
  OAI22X1 reg_in_U355 ( .A0(reg_in_n926), .A1(reg_in_n90), .B0(reg_in_n10), 
        .B1(reg_in_n927), .Y(reg_in_n621) );
  OAI22X1 reg_in_U354 ( .A0(reg_in_n927), .A1(reg_in_n91), .B0(reg_in_n10), 
        .B1(reg_in_n928), .Y(reg_in_n620) );
  OAI22X1 reg_in_U353 ( .A0(reg_in_n928), .A1(reg_in_n91), .B0(reg_in_n10), 
        .B1(reg_in_n929), .Y(reg_in_n619) );
  OAI22X1 reg_in_U352 ( .A0(reg_in_n929), .A1(reg_in_n92), .B0(reg_in_n10), 
        .B1(reg_in_n930), .Y(reg_in_n618) );
  OAI22X1 reg_in_U351 ( .A0(reg_in_n930), .A1(reg_in_n92), .B0(reg_in_n10), 
        .B1(reg_in_n931), .Y(reg_in_n617) );
  OAI22X1 reg_in_U350 ( .A0(reg_in_n931), .A1(reg_in_n93), .B0(reg_in_n10), 
        .B1(reg_in_n932), .Y(reg_in_n616) );
  OAI22X1 reg_in_U349 ( .A0(reg_in_n932), .A1(reg_in_n93), .B0(reg_in_n10), 
        .B1(reg_in_n933), .Y(reg_in_n615) );
  OAI22X1 reg_in_U348 ( .A0(reg_in_n933), .A1(reg_in_n94), .B0(reg_in_n10), 
        .B1(reg_in_n934), .Y(reg_in_n614) );
  OAI22X1 reg_in_U347 ( .A0(reg_in_n934), .A1(reg_in_n94), .B0(reg_in_n10), 
        .B1(reg_in_n935), .Y(reg_in_n613) );
  OAI22X1 reg_in_U346 ( .A0(reg_in_n937), .A1(reg_in_n94), .B0(reg_in_n10), 
        .B1(reg_in_n938), .Y(reg_in_n610) );
  OAI22X1 reg_in_U345 ( .A0(reg_in_n938), .A1(reg_in_n95), .B0(reg_in_n9), 
        .B1(reg_in_n939), .Y(reg_in_n609) );
  OAI22X1 reg_in_U344 ( .A0(reg_in_n939), .A1(reg_in_n95), .B0(reg_in_n9), 
        .B1(reg_in_n940), .Y(reg_in_n608) );
  OAI22X1 reg_in_U343 ( .A0(reg_in_n940), .A1(reg_in_n96), .B0(reg_in_n9), 
        .B1(reg_in_n941), .Y(reg_in_n607) );
  OAI22X1 reg_in_U342 ( .A0(reg_in_n941), .A1(reg_in_n96), .B0(reg_in_n9), 
        .B1(reg_in_n942), .Y(reg_in_n606) );
  OAI22X1 reg_in_U341 ( .A0(reg_in_n942), .A1(reg_in_n97), .B0(reg_in_n9), 
        .B1(reg_in_n943), .Y(reg_in_n605) );
  OAI22X1 reg_in_U340 ( .A0(reg_in_n943), .A1(reg_in_n97), .B0(reg_in_n9), 
        .B1(reg_in_n944), .Y(reg_in_n604) );
  OAI22X1 reg_in_U339 ( .A0(reg_in_n944), .A1(reg_in_n98), .B0(reg_in_n9), 
        .B1(reg_in_n945), .Y(reg_in_n603) );
  OAI22X1 reg_in_U338 ( .A0(reg_in_n945), .A1(reg_in_n98), .B0(reg_in_n9), 
        .B1(reg_in_n946), .Y(reg_in_n602) );
  OAI22X1 reg_in_U337 ( .A0(reg_in_n946), .A1(reg_in_n99), .B0(reg_in_n9), 
        .B1(reg_in_n947), .Y(reg_in_n601) );
  OAI22X1 reg_in_U336 ( .A0(reg_in_n947), .A1(reg_in_n99), .B0(reg_in_n9), 
        .B1(reg_in_n948), .Y(reg_in_n600) );
  OAI22X1 reg_in_U335 ( .A0(reg_in_n948), .A1(reg_in_n100), .B0(reg_in_n9), 
        .B1(reg_in_n949), .Y(reg_in_n599) );
  OAI22X1 reg_in_U334 ( .A0(reg_in_n949), .A1(reg_in_n100), .B0(reg_in_n9), 
        .B1(reg_in_n950), .Y(reg_in_n598) );
  OAI22X1 reg_in_U333 ( .A0(reg_in_n950), .A1(reg_in_n101), .B0(reg_in_n9), 
        .B1(reg_in_n951), .Y(reg_in_n597) );
  OAI22X1 reg_in_U332 ( .A0(reg_in_n951), .A1(reg_in_n101), .B0(reg_in_n8), 
        .B1(reg_in_n952), .Y(reg_in_n596) );
  OAI22X1 reg_in_U331 ( .A0(reg_in_n952), .A1(reg_in_n102), .B0(reg_in_n8), 
        .B1(reg_in_n953), .Y(reg_in_n595) );
  OAI22X1 reg_in_U330 ( .A0(reg_in_n953), .A1(reg_in_n102), .B0(reg_in_n8), 
        .B1(reg_in_n954), .Y(reg_in_n594) );
  OAI22X1 reg_in_U329 ( .A0(reg_in_n954), .A1(reg_in_n103), .B0(reg_in_n8), 
        .B1(reg_in_n955), .Y(reg_in_n593) );
  OAI22X1 reg_in_U328 ( .A0(reg_in_n955), .A1(reg_in_n103), .B0(reg_in_n8), 
        .B1(reg_in_n956), .Y(reg_in_n592) );
  OAI22X1 reg_in_U327 ( .A0(reg_in_n956), .A1(reg_in_n104), .B0(reg_in_n8), 
        .B1(reg_in_n957), .Y(reg_in_n591) );
  OAI22X1 reg_in_U326 ( .A0(reg_in_n957), .A1(reg_in_n104), .B0(reg_in_n8), 
        .B1(reg_in_n958), .Y(reg_in_n590) );
  OAI22X1 reg_in_U325 ( .A0(reg_in_n958), .A1(reg_in_n105), .B0(reg_in_n8), 
        .B1(reg_in_n959), .Y(reg_in_n589) );
  OAI22X1 reg_in_U324 ( .A0(reg_in_n959), .A1(reg_in_n105), .B0(reg_in_n8), 
        .B1(reg_in_n960), .Y(reg_in_n588) );
  OAI22X1 reg_in_U323 ( .A0(reg_in_n960), .A1(reg_in_n106), .B0(reg_in_n8), 
        .B1(reg_in_n961), .Y(reg_in_n587) );
  OAI22X1 reg_in_U322 ( .A0(reg_in_n961), .A1(reg_in_n106), .B0(reg_in_n8), 
        .B1(reg_in_n962), .Y(reg_in_n586) );
  OAI22X1 reg_in_U321 ( .A0(reg_in_n962), .A1(reg_in_n107), .B0(reg_in_n8), 
        .B1(reg_in_n963), .Y(reg_in_n585) );
  OAI22X1 reg_in_U320 ( .A0(reg_in_n963), .A1(reg_in_n107), .B0(reg_in_n8), 
        .B1(reg_in_n964), .Y(reg_in_n584) );
  OAI22X1 reg_in_U319 ( .A0(reg_in_n964), .A1(reg_in_n108), .B0(reg_in_n7), 
        .B1(reg_in_n965), .Y(reg_in_n583) );
  OAI22X1 reg_in_U318 ( .A0(reg_in_n965), .A1(reg_in_n108), .B0(reg_in_n7), 
        .B1(reg_in_n966), .Y(reg_in_n582) );
  OAI22X1 reg_in_U317 ( .A0(reg_in_n966), .A1(reg_in_n108), .B0(reg_in_n7), 
        .B1(reg_in_n967), .Y(reg_in_n581) );
  OAI22X1 reg_in_U316 ( .A0(reg_in_n969), .A1(reg_in_n109), .B0(reg_in_n7), 
        .B1(reg_in_n970), .Y(reg_in_n578) );
  OAI22X1 reg_in_U315 ( .A0(reg_in_n970), .A1(reg_in_n109), .B0(reg_in_n15), 
        .B1(reg_in_n971), .Y(reg_in_n577) );
  OAI22X1 reg_in_U314 ( .A0(reg_in_n971), .A1(reg_in_n110), .B0(reg_in_n7), 
        .B1(reg_in_n972), .Y(reg_in_n576) );
  OAI22X1 reg_in_U313 ( .A0(reg_in_n972), .A1(reg_in_n110), .B0(reg_in_n7), 
        .B1(reg_in_n973), .Y(reg_in_n575) );
  OAI22X1 reg_in_U312 ( .A0(reg_in_n973), .A1(reg_in_n111), .B0(reg_in_n7), 
        .B1(reg_in_n974), .Y(reg_in_n574) );
  OAI22X1 reg_in_U311 ( .A0(reg_in_n974), .A1(reg_in_n111), .B0(reg_in_n7), 
        .B1(reg_in_n975), .Y(reg_in_n573) );
  OAI22X1 reg_in_U310 ( .A0(reg_in_n975), .A1(reg_in_n112), .B0(reg_in_n6), 
        .B1(reg_in_n976), .Y(reg_in_n572) );
  OAI22X1 reg_in_U309 ( .A0(reg_in_n976), .A1(reg_in_n112), .B0(reg_in_n6), 
        .B1(reg_in_n977), .Y(reg_in_n571) );
  OAI22X1 reg_in_U308 ( .A0(reg_in_n977), .A1(reg_in_n113), .B0(reg_in_n6), 
        .B1(reg_in_n978), .Y(reg_in_n570) );
  OAI22X1 reg_in_U307 ( .A0(reg_in_n978), .A1(reg_in_n113), .B0(reg_in_n6), 
        .B1(reg_in_n979), .Y(reg_in_n569) );
  OAI22X1 reg_in_U306 ( .A0(reg_in_n979), .A1(reg_in_n114), .B0(reg_in_n6), 
        .B1(reg_in_n980), .Y(reg_in_n568) );
  OAI22X1 reg_in_U305 ( .A0(reg_in_n980), .A1(reg_in_n114), .B0(reg_in_n6), 
        .B1(reg_in_n981), .Y(reg_in_n567) );
  OAI22X1 reg_in_U304 ( .A0(reg_in_n981), .A1(reg_in_n115), .B0(reg_in_n6), 
        .B1(reg_in_n982), .Y(reg_in_n566) );
  OAI22X1 reg_in_U303 ( .A0(reg_in_n982), .A1(reg_in_n115), .B0(reg_in_n6), 
        .B1(reg_in_n983), .Y(reg_in_n565) );
  OAI22X1 reg_in_U302 ( .A0(reg_in_n983), .A1(reg_in_n116), .B0(reg_in_n6), 
        .B1(reg_in_n984), .Y(reg_in_n564) );
  OAI22X1 reg_in_U301 ( .A0(reg_in_n984), .A1(reg_in_n116), .B0(reg_in_n6), 
        .B1(reg_in_n985), .Y(reg_in_n563) );
  OAI22X1 reg_in_U300 ( .A0(reg_in_n985), .A1(reg_in_n117), .B0(reg_in_n6), 
        .B1(reg_in_n986), .Y(reg_in_n562) );
  OAI22X1 reg_in_U299 ( .A0(reg_in_n986), .A1(reg_in_n117), .B0(reg_in_n6), 
        .B1(reg_in_n987), .Y(reg_in_n561) );
  OAI22X1 reg_in_U298 ( .A0(reg_in_n987), .A1(reg_in_n118), .B0(reg_in_n6), 
        .B1(reg_in_n988), .Y(reg_in_n560) );
  OAI22X1 reg_in_U297 ( .A0(reg_in_n988), .A1(reg_in_n118), .B0(reg_in_n5), 
        .B1(reg_in_n989), .Y(reg_in_n559) );
  OAI22X1 reg_in_U296 ( .A0(reg_in_n989), .A1(reg_in_n119), .B0(reg_in_n5), 
        .B1(reg_in_n990), .Y(reg_in_n558) );
  OAI22X1 reg_in_U295 ( .A0(reg_in_n990), .A1(reg_in_n119), .B0(reg_in_n5), 
        .B1(reg_in_n991), .Y(reg_in_n557) );
  OAI22X1 reg_in_U294 ( .A0(reg_in_n991), .A1(reg_in_n120), .B0(reg_in_n5), 
        .B1(reg_in_n992), .Y(reg_in_n556) );
  OAI22X1 reg_in_U293 ( .A0(reg_in_n992), .A1(reg_in_n120), .B0(reg_in_n5), 
        .B1(reg_in_n993), .Y(reg_in_n555) );
  OAI22X1 reg_in_U292 ( .A0(reg_in_n993), .A1(reg_in_n121), .B0(reg_in_n5), 
        .B1(reg_in_n994), .Y(reg_in_n554) );
  OAI22X1 reg_in_U291 ( .A0(reg_in_n994), .A1(reg_in_n121), .B0(reg_in_n5), 
        .B1(reg_in_n995), .Y(reg_in_n553) );
  OAI22X1 reg_in_U290 ( .A0(reg_in_n995), .A1(reg_in_n122), .B0(reg_in_n5), 
        .B1(reg_in_n996), .Y(reg_in_n552) );
  OAI22X1 reg_in_U289 ( .A0(reg_in_n996), .A1(reg_in_n122), .B0(reg_in_n5), 
        .B1(reg_in_n997), .Y(reg_in_n551) );
  OAI22X1 reg_in_U288 ( .A0(reg_in_n997), .A1(reg_in_n123), .B0(reg_in_n5), 
        .B1(reg_in_n998), .Y(reg_in_n550) );
  OAI22X1 reg_in_U287 ( .A0(reg_in_n998), .A1(reg_in_n123), .B0(reg_in_n5), 
        .B1(reg_in_n999), .Y(reg_in_n549) );
  OAI22X1 reg_in_U286 ( .A0(reg_in_n1001), .A1(reg_in_n124), .B0(reg_in_n4), 
        .B1(reg_in_n1002), .Y(reg_in_n546) );
  OAI22X1 reg_in_U285 ( .A0(reg_in_n1002), .A1(reg_in_n125), .B0(reg_in_n4), 
        .B1(reg_in_n1003), .Y(reg_in_n545) );
  OAI22X1 reg_in_U284 ( .A0(reg_in_n1003), .A1(reg_in_n125), .B0(reg_in_n4), 
        .B1(reg_in_n1004), .Y(reg_in_n544) );
  OAI22X1 reg_in_U283 ( .A0(reg_in_n1004), .A1(reg_in_n126), .B0(reg_in_n4), 
        .B1(reg_in_n1005), .Y(reg_in_n543) );
  OAI22X1 reg_in_U282 ( .A0(reg_in_n1005), .A1(reg_in_n126), .B0(reg_in_n4), 
        .B1(reg_in_n1006), .Y(reg_in_n542) );
  OAI22X1 reg_in_U281 ( .A0(reg_in_n1006), .A1(reg_in_n127), .B0(reg_in_n4), 
        .B1(reg_in_n1007), .Y(reg_in_n541) );
  OAI22X1 reg_in_U280 ( .A0(reg_in_n1007), .A1(reg_in_n127), .B0(reg_in_n4), 
        .B1(reg_in_n1008), .Y(reg_in_n540) );
  OAI22X1 reg_in_U279 ( .A0(reg_in_n1008), .A1(reg_in_n128), .B0(reg_in_n4), 
        .B1(reg_in_n1009), .Y(reg_in_n539) );
  OAI22X1 reg_in_U278 ( .A0(reg_in_n1009), .A1(reg_in_n128), .B0(reg_in_n4), 
        .B1(reg_in_n1010), .Y(reg_in_n538) );
  OAI22X1 reg_in_U277 ( .A0(reg_in_n1010), .A1(reg_in_n129), .B0(reg_in_n4), 
        .B1(reg_in_n1011), .Y(reg_in_n537) );
  OAI22X1 reg_in_U276 ( .A0(reg_in_n1011), .A1(reg_in_n129), .B0(reg_in_n4), 
        .B1(reg_in_n1012), .Y(reg_in_n536) );
  OAI22X1 reg_in_U275 ( .A0(reg_in_n1012), .A1(reg_in_n130), .B0(reg_in_n4), 
        .B1(reg_in_n1013), .Y(reg_in_n535) );
  OAI22X1 reg_in_U274 ( .A0(reg_in_n1013), .A1(reg_in_n130), .B0(reg_in_n4), 
        .B1(reg_in_n1014), .Y(reg_in_n534) );
  OAI22X1 reg_in_U273 ( .A0(reg_in_n1014), .A1(reg_in_n131), .B0(reg_in_n3), 
        .B1(reg_in_n1015), .Y(reg_in_n533) );
  OAI22X1 reg_in_U272 ( .A0(reg_in_n1015), .A1(reg_in_n131), .B0(reg_in_n3), 
        .B1(reg_in_n1016), .Y(reg_in_n532) );
  OAI22X1 reg_in_U271 ( .A0(reg_in_n1016), .A1(reg_in_n132), .B0(reg_in_n3), 
        .B1(reg_in_n1017), .Y(reg_in_n531) );
  OAI22X1 reg_in_U270 ( .A0(reg_in_n1017), .A1(reg_in_n132), .B0(reg_in_n3), 
        .B1(reg_in_n1018), .Y(reg_in_n530) );
  OAI22X1 reg_in_U269 ( .A0(reg_in_n1018), .A1(reg_in_n133), .B0(reg_in_n3), 
        .B1(reg_in_n1019), .Y(reg_in_n529) );
  OAI22X1 reg_in_U268 ( .A0(reg_in_n1019), .A1(reg_in_n133), .B0(reg_in_n3), 
        .B1(reg_in_n1020), .Y(reg_in_n528) );
  OAI22X1 reg_in_U267 ( .A0(reg_in_n1020), .A1(reg_in_n134), .B0(reg_in_n3), 
        .B1(reg_in_n1021), .Y(reg_in_n527) );
  OAI22X1 reg_in_U266 ( .A0(reg_in_n1021), .A1(reg_in_n134), .B0(reg_in_n3), 
        .B1(reg_in_n1022), .Y(reg_in_n526) );
  OAI22X1 reg_in_U265 ( .A0(reg_in_n1022), .A1(reg_in_n135), .B0(reg_in_n3), 
        .B1(reg_in_n1023), .Y(reg_in_n525) );
  OAI22X1 reg_in_U264 ( .A0(reg_in_n1023), .A1(reg_in_n135), .B0(reg_in_n2), 
        .B1(reg_in_n1024), .Y(reg_in_n524) );
  OAI22X1 reg_in_U263 ( .A0(reg_in_n1024), .A1(reg_in_n136), .B0(reg_in_n5), 
        .B1(reg_in_n1025), .Y(reg_in_n523) );
  OAI22X1 reg_in_U262 ( .A0(reg_in_n1025), .A1(reg_in_n136), .B0(reg_in_n7), 
        .B1(reg_in_n1026), .Y(reg_in_n522) );
  OAI22X1 reg_in_U261 ( .A0(reg_in_n1026), .A1(reg_in_n137), .B0(reg_in_n10), 
        .B1(reg_in_n1027), .Y(reg_in_n521) );
  OAI22X1 reg_in_U260 ( .A0(reg_in_n1027), .A1(reg_in_n137), .B0(reg_in_n12), 
        .B1(reg_in_n1028), .Y(reg_in_n520) );
  OAI22X1 reg_in_U259 ( .A0(reg_in_n1028), .A1(reg_in_n138), .B0(reg_in_n15), 
        .B1(reg_in_n1029), .Y(reg_in_n519) );
  OAI22X1 reg_in_U258 ( .A0(reg_in_n1029), .A1(reg_in_n138), .B0(reg_in_n12), 
        .B1(reg_in_n1030), .Y(reg_in_n518) );
  OAI22X1 reg_in_U257 ( .A0(reg_in_n1030), .A1(reg_in_n117), .B0(reg_in_n12), 
        .B1(reg_in_n1031), .Y(reg_in_n517) );
  INVX1 reg_in_U256 ( .A(reg_in_n211), .Y(reg_in_n188) );
  INVX1 reg_in_U255 ( .A(reg_in_n216), .Y(reg_in_n189) );
  INVX1 reg_in_U254 ( .A(reg_in_n216), .Y(reg_in_n190) );
  INVX1 reg_in_U253 ( .A(reg_in_n216), .Y(reg_in_n191) );
  INVX1 reg_in_U252 ( .A(reg_in_n215), .Y(reg_in_n192) );
  INVX1 reg_in_U251 ( .A(reg_in_n215), .Y(reg_in_n193) );
  INVX1 reg_in_U250 ( .A(reg_in_n215), .Y(reg_in_n194) );
  INVX1 reg_in_U249 ( .A(reg_in_n214), .Y(reg_in_n195) );
  INVX1 reg_in_U248 ( .A(reg_in_n214), .Y(reg_in_n196) );
  INVX1 reg_in_U247 ( .A(reg_in_n214), .Y(reg_in_n197) );
  INVX1 reg_in_U246 ( .A(reg_in_n213), .Y(reg_in_n198) );
  INVX1 reg_in_U245 ( .A(reg_in_n213), .Y(reg_in_n199) );
  INVX1 reg_in_U244 ( .A(reg_in_n213), .Y(reg_in_n200) );
  INVX1 reg_in_U243 ( .A(reg_in_n212), .Y(reg_in_n201) );
  INVX1 reg_in_U242 ( .A(reg_in_n212), .Y(reg_in_n202) );
  INVX1 reg_in_U241 ( .A(reg_in_n212), .Y(reg_in_n203) );
  INVX1 reg_in_U240 ( .A(reg_in_n211), .Y(reg_in_n204) );
  INVX1 reg_in_U239 ( .A(reg_in_n211), .Y(reg_in_n205) );
  INVX1 reg_in_U238 ( .A(reg_in_n211), .Y(reg_in_n206) );
  INVX1 reg_in_U237 ( .A(reg_in_n210), .Y(reg_in_n207) );
  INVX1 reg_in_U236 ( .A(reg_in_n210), .Y(reg_in_n208) );
  INVX1 reg_in_U235 ( .A(reg_in_n219), .Y(reg_in_n218) );
  INVX1 reg_in_U234 ( .A(reg_in_n219), .Y(reg_in_n217) );
  INVX1 reg_in_U233 ( .A(reg_in_n210), .Y(reg_in_n209) );
  INVX1 reg_in_U232 ( .A(reg_in_n209), .Y(reg_in_n149) );
  INVX1 reg_in_U231 ( .A(reg_in_n149), .Y(reg_in_n148) );
  INVX1 reg_in_U230 ( .A(reg_in_n149), .Y(reg_in_n147) );
  INVX1 reg_in_U229 ( .A(reg_in_n218), .Y(reg_in_n776) );
  INVX1 reg_in_U228 ( .A(reg_in_n217), .Y(reg_in_n257) );
  INVX1 reg_in_U227 ( .A(reg_in_n218), .Y(reg_in_n773) );
  INVX1 reg_in_U226 ( .A(reg_in_n218), .Y(reg_in_n774) );
  INVX1 reg_in_U225 ( .A(reg_in_n217), .Y(reg_in_n254) );
  INVX1 reg_in_U224 ( .A(reg_in_n218), .Y(reg_in_n775) );
  INVX1 reg_in_U223 ( .A(reg_in_n217), .Y(reg_in_n255) );
  INVX1 reg_in_U222 ( .A(reg_in_n217), .Y(reg_in_n256) );
  INVX1 reg_in_U221 ( .A(reg_in_n217), .Y(reg_in_n259) );
  INVX1 reg_in_U220 ( .A(reg_in_n218), .Y(reg_in_n772) );
  INVX1 reg_in_U219 ( .A(reg_in_n188), .Y(reg_in_n187) );
  INVX1 reg_in_U218 ( .A(reg_in_n188), .Y(reg_in_n186) );
  INVX1 reg_in_U217 ( .A(reg_in_n188), .Y(reg_in_n185) );
  INVX1 reg_in_U216 ( .A(reg_in_n188), .Y(reg_in_n184) );
  INVX1 reg_in_U215 ( .A(reg_in_n189), .Y(reg_in_n183) );
  INVX1 reg_in_U214 ( .A(reg_in_n190), .Y(reg_in_n182) );
  INVX1 reg_in_U213 ( .A(reg_in_n191), .Y(reg_in_n181) );
  INVX1 reg_in_U212 ( .A(reg_in_n191), .Y(reg_in_n180) );
  INVX1 reg_in_U211 ( .A(reg_in_n192), .Y(reg_in_n179) );
  INVX1 reg_in_U210 ( .A(reg_in_n192), .Y(reg_in_n178) );
  INVX1 reg_in_U209 ( .A(reg_in_n193), .Y(reg_in_n177) );
  INVX1 reg_in_U208 ( .A(reg_in_n193), .Y(reg_in_n176) );
  INVX1 reg_in_U207 ( .A(reg_in_n194), .Y(reg_in_n175) );
  INVX1 reg_in_U206 ( .A(reg_in_n195), .Y(reg_in_n174) );
  INVX1 reg_in_U205 ( .A(reg_in_n195), .Y(reg_in_n173) );
  INVX1 reg_in_U204 ( .A(reg_in_n196), .Y(reg_in_n172) );
  INVX1 reg_in_U203 ( .A(reg_in_n196), .Y(reg_in_n171) );
  INVX1 reg_in_U202 ( .A(reg_in_n197), .Y(reg_in_n170) );
  INVX1 reg_in_U201 ( .A(reg_in_n198), .Y(reg_in_n169) );
  INVX1 reg_in_U200 ( .A(reg_in_n198), .Y(reg_in_n168) );
  INVX1 reg_in_U199 ( .A(reg_in_n199), .Y(reg_in_n167) );
  INVX1 reg_in_U198 ( .A(reg_in_n200), .Y(reg_in_n166) );
  INVX1 reg_in_U197 ( .A(reg_in_n200), .Y(reg_in_n165) );
  INVX1 reg_in_U196 ( .A(reg_in_n201), .Y(reg_in_n164) );
  INVX1 reg_in_U195 ( .A(reg_in_n201), .Y(reg_in_n163) );
  INVX1 reg_in_U194 ( .A(reg_in_n202), .Y(reg_in_n162) );
  INVX1 reg_in_U193 ( .A(reg_in_n203), .Y(reg_in_n161) );
  INVX1 reg_in_U192 ( .A(reg_in_n203), .Y(reg_in_n160) );
  INVX1 reg_in_U191 ( .A(reg_in_n204), .Y(reg_in_n159) );
  INVX1 reg_in_U190 ( .A(reg_in_n204), .Y(reg_in_n158) );
  INVX1 reg_in_U189 ( .A(reg_in_n205), .Y(reg_in_n157) );
  INVX1 reg_in_U188 ( .A(reg_in_n205), .Y(reg_in_n156) );
  INVX1 reg_in_U187 ( .A(reg_in_n206), .Y(reg_in_n155) );
  INVX1 reg_in_U186 ( .A(reg_in_n206), .Y(reg_in_n154) );
  INVX1 reg_in_U185 ( .A(reg_in_n207), .Y(reg_in_n153) );
  INVX1 reg_in_U184 ( .A(reg_in_n207), .Y(reg_in_n152) );
  INVX1 reg_in_U183 ( .A(reg_in_n208), .Y(reg_in_n151) );
  INVX1 reg_in_U182 ( .A(reg_in_n208), .Y(reg_in_n150) );
  INVX1 reg_in_U181 ( .A(reg_in_n152), .Y(reg_in_n139) );
  INVX1 reg_in_U180 ( .A(reg_in_n151), .Y(reg_in_n141) );
  INVX1 reg_in_U179 ( .A(reg_in_n150), .Y(reg_in_n146) );
  INVX1 reg_in_U178 ( .A(reg_in_n150), .Y(reg_in_n144) );
  INVX1 reg_in_U177 ( .A(reg_in_n150), .Y(reg_in_n145) );
  INVX1 reg_in_U176 ( .A(reg_in_n151), .Y(reg_in_n143) );
  INVX1 reg_in_U175 ( .A(reg_in_n151), .Y(reg_in_n142) );
  INVX1 reg_in_U174 ( .A(reg_in_n152), .Y(reg_in_n140) );
  INVX1 reg_in_U173 ( .A(reg_in_n187), .Y(reg_in_n22) );
  INVX1 reg_in_U172 ( .A(reg_in_n187), .Y(reg_in_n23) );
  INVX1 reg_in_U171 ( .A(reg_in_n187), .Y(reg_in_n24) );
  INVX1 reg_in_U170 ( .A(reg_in_n186), .Y(reg_in_n25) );
  INVX1 reg_in_U169 ( .A(reg_in_n186), .Y(reg_in_n26) );
  INVX1 reg_in_U168 ( .A(reg_in_n186), .Y(reg_in_n27) );
  INVX1 reg_in_U167 ( .A(reg_in_n185), .Y(reg_in_n28) );
  INVX1 reg_in_U166 ( .A(reg_in_n185), .Y(reg_in_n29) );
  INVX1 reg_in_U165 ( .A(reg_in_n185), .Y(reg_in_n30) );
  INVX1 reg_in_U164 ( .A(reg_in_n184), .Y(reg_in_n31) );
  INVX1 reg_in_U163 ( .A(reg_in_n184), .Y(reg_in_n32) );
  INVX1 reg_in_U162 ( .A(reg_in_n184), .Y(reg_in_n33) );
  INVX1 reg_in_U161 ( .A(reg_in_n183), .Y(reg_in_n34) );
  INVX1 reg_in_U160 ( .A(reg_in_n183), .Y(reg_in_n35) );
  INVX1 reg_in_U159 ( .A(reg_in_n183), .Y(reg_in_n36) );
  INVX1 reg_in_U158 ( .A(reg_in_n183), .Y(reg_in_n37) );
  INVX1 reg_in_U157 ( .A(reg_in_n183), .Y(reg_in_n38) );
  INVX1 reg_in_U156 ( .A(reg_in_n182), .Y(reg_in_n39) );
  INVX1 reg_in_U155 ( .A(reg_in_n182), .Y(reg_in_n40) );
  INVX1 reg_in_U154 ( .A(reg_in_n182), .Y(reg_in_n41) );
  INVX1 reg_in_U153 ( .A(reg_in_n182), .Y(reg_in_n42) );
  INVX1 reg_in_U152 ( .A(reg_in_n182), .Y(reg_in_n43) );
  INVX1 reg_in_U151 ( .A(reg_in_n181), .Y(reg_in_n44) );
  INVX1 reg_in_U150 ( .A(reg_in_n181), .Y(reg_in_n45) );
  INVX1 reg_in_U149 ( .A(reg_in_n181), .Y(reg_in_n46) );
  INVX1 reg_in_U148 ( .A(reg_in_n180), .Y(reg_in_n47) );
  INVX1 reg_in_U147 ( .A(reg_in_n180), .Y(reg_in_n48) );
  INVX1 reg_in_U146 ( .A(reg_in_n180), .Y(reg_in_n49) );
  INVX1 reg_in_U145 ( .A(reg_in_n179), .Y(reg_in_n50) );
  INVX1 reg_in_U144 ( .A(reg_in_n179), .Y(reg_in_n51) );
  INVX1 reg_in_U143 ( .A(reg_in_n179), .Y(reg_in_n52) );
  INVX1 reg_in_U142 ( .A(reg_in_n178), .Y(reg_in_n53) );
  INVX1 reg_in_U141 ( .A(reg_in_n178), .Y(reg_in_n54) );
  INVX1 reg_in_U140 ( .A(reg_in_n178), .Y(reg_in_n55) );
  INVX1 reg_in_U139 ( .A(reg_in_n177), .Y(reg_in_n56) );
  INVX1 reg_in_U138 ( .A(reg_in_n177), .Y(reg_in_n57) );
  INVX1 reg_in_U137 ( .A(reg_in_n177), .Y(reg_in_n58) );
  INVX1 reg_in_U136 ( .A(reg_in_n176), .Y(reg_in_n59) );
  INVX1 reg_in_U135 ( .A(reg_in_n176), .Y(reg_in_n60) );
  INVX1 reg_in_U134 ( .A(reg_in_n176), .Y(reg_in_n61) );
  INVX1 reg_in_U133 ( .A(reg_in_n175), .Y(reg_in_n62) );
  INVX1 reg_in_U132 ( .A(reg_in_n175), .Y(reg_in_n63) );
  INVX1 reg_in_U131 ( .A(reg_in_n175), .Y(reg_in_n64) );
  INVX1 reg_in_U130 ( .A(reg_in_n175), .Y(reg_in_n65) );
  INVX1 reg_in_U129 ( .A(reg_in_n175), .Y(reg_in_n66) );
  INVX1 reg_in_U128 ( .A(reg_in_n174), .Y(reg_in_n67) );
  INVX1 reg_in_U127 ( .A(reg_in_n174), .Y(reg_in_n68) );
  INVX1 reg_in_U126 ( .A(reg_in_n174), .Y(reg_in_n69) );
  INVX1 reg_in_U125 ( .A(reg_in_n173), .Y(reg_in_n70) );
  INVX1 reg_in_U124 ( .A(reg_in_n173), .Y(reg_in_n71) );
  INVX1 reg_in_U123 ( .A(reg_in_n173), .Y(reg_in_n72) );
  INVX1 reg_in_U122 ( .A(reg_in_n172), .Y(reg_in_n73) );
  INVX1 reg_in_U121 ( .A(reg_in_n172), .Y(reg_in_n74) );
  INVX1 reg_in_U120 ( .A(reg_in_n172), .Y(reg_in_n75) );
  INVX1 reg_in_U119 ( .A(reg_in_n171), .Y(reg_in_n76) );
  INVX1 reg_in_U118 ( .A(reg_in_n171), .Y(reg_in_n77) );
  INVX1 reg_in_U117 ( .A(reg_in_n171), .Y(reg_in_n78) );
  INVX1 reg_in_U116 ( .A(reg_in_n170), .Y(reg_in_n79) );
  INVX1 reg_in_U115 ( .A(reg_in_n170), .Y(reg_in_n80) );
  INVX1 reg_in_U114 ( .A(reg_in_n170), .Y(reg_in_n81) );
  INVX1 reg_in_U113 ( .A(reg_in_n170), .Y(reg_in_n82) );
  INVX1 reg_in_U112 ( .A(reg_in_n170), .Y(reg_in_n83) );
  INVX1 reg_in_U111 ( .A(reg_in_n169), .Y(reg_in_n84) );
  INVX1 reg_in_U110 ( .A(reg_in_n169), .Y(reg_in_n85) );
  INVX1 reg_in_U109 ( .A(reg_in_n169), .Y(reg_in_n86) );
  INVX1 reg_in_U108 ( .A(reg_in_n168), .Y(reg_in_n87) );
  INVX1 reg_in_U107 ( .A(reg_in_n168), .Y(reg_in_n88) );
  INVX1 reg_in_U106 ( .A(reg_in_n168), .Y(reg_in_n89) );
  INVX1 reg_in_U105 ( .A(reg_in_n167), .Y(reg_in_n90) );
  INVX1 reg_in_U104 ( .A(reg_in_n167), .Y(reg_in_n91) );
  INVX1 reg_in_U103 ( .A(reg_in_n167), .Y(reg_in_n92) );
  INVX1 reg_in_U102 ( .A(reg_in_n167), .Y(reg_in_n93) );
  INVX1 reg_in_U101 ( .A(reg_in_n167), .Y(reg_in_n94) );
  INVX1 reg_in_U100 ( .A(reg_in_n166), .Y(reg_in_n95) );
  INVX1 reg_in_U99 ( .A(reg_in_n166), .Y(reg_in_n96) );
  INVX1 reg_in_U98 ( .A(reg_in_n166), .Y(reg_in_n97) );
  INVX1 reg_in_U97 ( .A(reg_in_n165), .Y(reg_in_n98) );
  INVX1 reg_in_U96 ( .A(reg_in_n165), .Y(reg_in_n99) );
  INVX1 reg_in_U95 ( .A(reg_in_n165), .Y(reg_in_n100) );
  INVX1 reg_in_U94 ( .A(reg_in_n164), .Y(reg_in_n101) );
  INVX1 reg_in_U93 ( .A(reg_in_n164), .Y(reg_in_n102) );
  INVX1 reg_in_U92 ( .A(reg_in_n164), .Y(reg_in_n103) );
  INVX1 reg_in_U91 ( .A(reg_in_n163), .Y(reg_in_n104) );
  INVX1 reg_in_U90 ( .A(reg_in_n163), .Y(reg_in_n105) );
  INVX1 reg_in_U89 ( .A(reg_in_n163), .Y(reg_in_n106) );
  INVX1 reg_in_U88 ( .A(reg_in_n162), .Y(reg_in_n107) );
  INVX1 reg_in_U87 ( .A(reg_in_n162), .Y(reg_in_n108) );
  INVX1 reg_in_U86 ( .A(reg_in_n162), .Y(reg_in_n109) );
  INVX1 reg_in_U85 ( .A(reg_in_n162), .Y(reg_in_n110) );
  INVX1 reg_in_U84 ( .A(reg_in_n162), .Y(reg_in_n111) );
  INVX1 reg_in_U83 ( .A(reg_in_n161), .Y(reg_in_n112) );
  INVX1 reg_in_U82 ( .A(reg_in_n161), .Y(reg_in_n113) );
  INVX1 reg_in_U81 ( .A(reg_in_n161), .Y(reg_in_n114) );
  INVX1 reg_in_U80 ( .A(reg_in_n160), .Y(reg_in_n115) );
  INVX1 reg_in_U79 ( .A(reg_in_n160), .Y(reg_in_n116) );
  INVX1 reg_in_U78 ( .A(reg_in_n160), .Y(reg_in_n117) );
  INVX1 reg_in_U77 ( .A(reg_in_n159), .Y(reg_in_n118) );
  INVX1 reg_in_U76 ( .A(reg_in_n159), .Y(reg_in_n119) );
  INVX1 reg_in_U75 ( .A(reg_in_n159), .Y(reg_in_n120) );
  INVX1 reg_in_U74 ( .A(reg_in_n158), .Y(reg_in_n121) );
  INVX1 reg_in_U73 ( .A(reg_in_n158), .Y(reg_in_n122) );
  INVX1 reg_in_U72 ( .A(reg_in_n158), .Y(reg_in_n123) );
  INVX1 reg_in_U71 ( .A(reg_in_n157), .Y(reg_in_n124) );
  INVX1 reg_in_U70 ( .A(reg_in_n157), .Y(reg_in_n125) );
  INVX1 reg_in_U69 ( .A(reg_in_n157), .Y(reg_in_n126) );
  INVX1 reg_in_U68 ( .A(reg_in_n156), .Y(reg_in_n127) );
  INVX1 reg_in_U67 ( .A(reg_in_n156), .Y(reg_in_n128) );
  INVX1 reg_in_U66 ( .A(reg_in_n156), .Y(reg_in_n129) );
  INVX1 reg_in_U65 ( .A(reg_in_n155), .Y(reg_in_n130) );
  INVX1 reg_in_U64 ( .A(reg_in_n155), .Y(reg_in_n131) );
  INVX1 reg_in_U63 ( .A(reg_in_n155), .Y(reg_in_n132) );
  INVX1 reg_in_U62 ( .A(reg_in_n154), .Y(reg_in_n133) );
  INVX1 reg_in_U61 ( .A(reg_in_n154), .Y(reg_in_n134) );
  INVX1 reg_in_U60 ( .A(reg_in_n154), .Y(reg_in_n135) );
  INVX1 reg_in_U59 ( .A(reg_in_n153), .Y(reg_in_n136) );
  INVX1 reg_in_U58 ( .A(reg_in_n153), .Y(reg_in_n137) );
  INVX1 reg_in_U57 ( .A(reg_in_n153), .Y(reg_in_n138) );
  INVX1 reg_in_U56 ( .A(reg_in_n257), .Y(reg_in_n253) );
  INVX1 reg_in_U55 ( .A(reg_in_n776), .Y(reg_in_n223) );
  INVX1 reg_in_U54 ( .A(reg_in_n776), .Y(reg_in_n220) );
  INVX1 reg_in_U53 ( .A(reg_in_n219), .Y(reg_in_n233) );
  INVX1 reg_in_U52 ( .A(reg_in_n219), .Y(reg_in_n232) );
  INVX1 reg_in_U51 ( .A(reg_in_n773), .Y(reg_in_n231) );
  INVX1 reg_in_U50 ( .A(reg_in_n774), .Y(reg_in_n230) );
  INVX1 reg_in_U49 ( .A(reg_in_n773), .Y(reg_in_n229) );
  INVX1 reg_in_U48 ( .A(reg_in_n773), .Y(reg_in_n228) );
  INVX1 reg_in_U47 ( .A(reg_in_n774), .Y(reg_in_n227) );
  INVX1 reg_in_U46 ( .A(reg_in_n774), .Y(reg_in_n226) );
  INVX1 reg_in_U45 ( .A(reg_in_n775), .Y(reg_in_n225) );
  INVX1 reg_in_U44 ( .A(reg_in_n775), .Y(reg_in_n224) );
  INVX1 reg_in_U43 ( .A(reg_in_n775), .Y(reg_in_n222) );
  INVX1 reg_in_U42 ( .A(reg_in_n776), .Y(reg_in_n221) );
  INVX1 reg_in_U41 ( .A(reg_in_n259), .Y(reg_in_n238) );
  INVX1 reg_in_U40 ( .A(reg_in_n259), .Y(reg_in_n239) );
  INVX1 reg_in_U39 ( .A(reg_in_n259), .Y(reg_in_n237) );
  INVX1 reg_in_U38 ( .A(reg_in_n772), .Y(reg_in_n236) );
  INVX1 reg_in_U37 ( .A(reg_in_n772), .Y(reg_in_n235) );
  INVX1 reg_in_U36 ( .A(reg_in_n772), .Y(reg_in_n234) );
  CLKINVX3 reg_in_U35 ( .A(reg_in_n148), .Y(reg_in_n21) );
  CLKINVX3 reg_in_U34 ( .A(reg_in_n254), .Y(reg_in_n240) );
  CLKINVX3 reg_in_U33 ( .A(reg_in_n255), .Y(reg_in_n241) );
  CLKINVX3 reg_in_U32 ( .A(reg_in_n257), .Y(reg_in_n242) );
  CLKINVX3 reg_in_U31 ( .A(reg_in_n256), .Y(reg_in_n243) );
  CLKINVX3 reg_in_U30 ( .A(reg_in_n257), .Y(reg_in_n244) );
  CLKINVX3 reg_in_U29 ( .A(reg_in_n257), .Y(reg_in_n245) );
  CLKINVX3 reg_in_U28 ( .A(reg_in_n256), .Y(reg_in_n252) );
  CLKINVX3 reg_in_U27 ( .A(reg_in_n254), .Y(reg_in_n251) );
  CLKINVX3 reg_in_U26 ( .A(reg_in_n254), .Y(reg_in_n250) );
  CLKINVX3 reg_in_U25 ( .A(reg_in_n255), .Y(reg_in_n249) );
  CLKINVX3 reg_in_U24 ( .A(reg_in_n255), .Y(reg_in_n248) );
  CLKINVX3 reg_in_U23 ( .A(reg_in_n256), .Y(reg_in_n247) );
  CLKINVX3 reg_in_U22 ( .A(reg_in_n256), .Y(reg_in_n246) );
  CLKINVX3 reg_in_U21 ( .A(reg_in_n148), .Y(reg_in_n20) );
  CLKINVX3 reg_in_U20 ( .A(reg_in_n147), .Y(reg_in_n19) );
  CLKINVX3 reg_in_U19 ( .A(reg_in_n147), .Y(reg_in_n18) );
  CLKINVX3 reg_in_U18 ( .A(reg_in_n141), .Y(reg_in_n7) );
  CLKINVX3 reg_in_U17 ( .A(reg_in_n146), .Y(reg_in_n17) );
  CLKINVX3 reg_in_U16 ( .A(reg_in_n139), .Y(reg_in_n3) );
  CLKINVX3 reg_in_U15 ( .A(reg_in_n144), .Y(reg_in_n12) );
  CLKINVX3 reg_in_U14 ( .A(reg_in_n144), .Y(reg_in_n13) );
  CLKINVX3 reg_in_U13 ( .A(reg_in_n146), .Y(reg_in_n16) );
  CLKINVX3 reg_in_U12 ( .A(reg_in_n145), .Y(reg_in_n15) );
  CLKINVX3 reg_in_U11 ( .A(reg_in_n145), .Y(reg_in_n14) );
  CLKINVX3 reg_in_U10 ( .A(reg_in_n143), .Y(reg_in_n11) );
  CLKINVX3 reg_in_U9 ( .A(reg_in_n143), .Y(reg_in_n10) );
  CLKINVX3 reg_in_U8 ( .A(reg_in_n142), .Y(reg_in_n9) );
  CLKINVX3 reg_in_U7 ( .A(reg_in_n142), .Y(reg_in_n8) );
  CLKINVX3 reg_in_U6 ( .A(reg_in_n141), .Y(reg_in_n6) );
  CLKINVX3 reg_in_U5 ( .A(reg_in_n140), .Y(reg_in_n5) );
  CLKINVX3 reg_in_U4 ( .A(reg_in_n140), .Y(reg_in_n4) );
  CLKINVX3 reg_in_U3 ( .A(reg_in_n139), .Y(reg_in_n2) );
  DFFRHQX1 reg_in_plain_key_out_reg_219_ ( .D(reg_in_n479), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[219]) );
  DFFRHQX1 reg_in_plain_key_out_reg_220_ ( .D(reg_in_n480), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[220]) );
  DFFRHQX1 reg_in_plain_key_out_reg_221_ ( .D(reg_in_n481), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[221]) );
  DFFRHQX1 reg_in_plain_key_out_reg_222_ ( .D(reg_in_n482), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[222]) );
  DFFRHQX1 reg_in_plain_key_out_reg_223_ ( .D(reg_in_n483), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[223]) );
  DFFRHQX1 reg_in_plain_key_out_reg_224_ ( .D(reg_in_n484), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[224]) );
  DFFRHQX1 reg_in_plain_key_out_reg_225_ ( .D(reg_in_n485), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[225]) );
  DFFRHQX1 reg_in_plain_key_out_reg_226_ ( .D(reg_in_n486), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[226]) );
  DFFRHQX1 reg_in_plain_key_out_reg_227_ ( .D(reg_in_n487), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[227]) );
  DFFRHQX1 reg_in_plain_key_out_reg_228_ ( .D(reg_in_n488), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[228]) );
  DFFRHQX1 reg_in_plain_key_out_reg_229_ ( .D(reg_in_n489), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[229]) );
  DFFRHQX1 reg_in_plain_key_out_reg_230_ ( .D(reg_in_n490), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[230]) );
  DFFRHQX1 reg_in_plain_key_out_reg_231_ ( .D(reg_in_n491), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[231]) );
  DFFRHQX1 reg_in_plain_key_out_reg_232_ ( .D(reg_in_n492), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[232]) );
  DFFRHQX1 reg_in_plain_key_out_reg_233_ ( .D(reg_in_n493), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[233]) );
  DFFRHQX1 reg_in_plain_key_out_reg_234_ ( .D(reg_in_n494), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[234]) );
  DFFRHQX1 reg_in_plain_key_out_reg_235_ ( .D(reg_in_n495), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[235]) );
  DFFRHQX1 reg_in_plain_key_out_reg_236_ ( .D(reg_in_n496), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[236]) );
  DFFRHQX1 reg_in_plain_key_out_reg_237_ ( .D(reg_in_n497), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[237]) );
  DFFRHQX1 reg_in_plain_key_out_reg_238_ ( .D(reg_in_n498), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[238]) );
  DFFRHQX1 reg_in_plain_key_out_reg_239_ ( .D(reg_in_n499), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[239]) );
  DFFRHQX1 reg_in_plain_key_out_reg_240_ ( .D(reg_in_n500), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[240]) );
  DFFRHQX1 reg_in_plain_key_out_reg_241_ ( .D(reg_in_n501), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[241]) );
  DFFRHQX1 reg_in_plain_key_out_reg_242_ ( .D(reg_in_n502), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[242]) );
  DFFRHQX1 reg_in_plain_key_out_reg_243_ ( .D(reg_in_n503), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[243]) );
  DFFRHQX1 reg_in_plain_key_out_reg_244_ ( .D(reg_in_n504), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[244]) );
  DFFRHQX1 reg_in_plain_key_out_reg_245_ ( .D(reg_in_n505), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[245]) );
  DFFRHQX1 reg_in_plain_key_out_reg_246_ ( .D(reg_in_n506), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[246]) );
  DFFRHQX1 reg_in_plain_key_out_reg_247_ ( .D(reg_in_n507), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[247]) );
  DFFRHQX1 reg_in_plain_key_out_reg_248_ ( .D(reg_in_n508), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[248]) );
  DFFRHQX1 reg_in_plain_key_out_reg_249_ ( .D(reg_in_n509), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[249]) );
  DFFRHQX1 reg_in_plain_key_out_reg_250_ ( .D(reg_in_n510), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[250]) );
  DFFRHQX1 reg_in_plain_key_out_reg_251_ ( .D(reg_in_n511), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[251]) );
  DFFRHQX1 reg_in_plain_key_out_reg_252_ ( .D(reg_in_n512), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[252]) );
  DFFRHQX1 reg_in_plain_key_out_reg_253_ ( .D(reg_in_n513), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[253]) );
  DFFRHQX1 reg_in_plain_key_out_reg_254_ ( .D(reg_in_n514), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[254]) );
  DFFRHQX1 reg_in_plain_key_out_reg_255_ ( .D(reg_in_n515), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[255]) );
  DFFRHQX1 reg_in_plain_key_out_reg_5_ ( .D(reg_in_n265), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[5]) );
  DFFRHQX1 reg_in_plain_key_out_reg_6_ ( .D(reg_in_n266), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[6]) );
  DFFRHQX1 reg_in_plain_key_out_reg_7_ ( .D(reg_in_n267), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[7]) );
  DFFRHQX1 reg_in_plain_key_out_reg_75_ ( .D(reg_in_n335), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[75]) );
  DFFRHQX1 reg_in_pbv1_reg ( .D(reg_in_pbv0), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(reg_in_pbv1) );
  DFFRHQX1 reg_in_pf1_reg ( .D(reg_in_pf0), .CK(clk_48Mhz), .RN(reset_n), .Q(
        reg_in_pf1) );
  DFFRHQX1 reg_in_pf0_reg ( .D(plain_finish), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(reg_in_pf0) );
  DFFRHQX1 reg_in_pbv0_reg ( .D(plain_byte_valid), .CK(clk_48Mhz), .RN(reset_n), .Q(reg_in_pbv0) );
  DFFRHQX1 reg_in_plain_key_out_reg_24_ ( .D(reg_in_n284), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[24]) );
  DFFRHQX1 reg_in_plain_key_out_reg_25_ ( .D(reg_in_n285), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[25]) );
  DFFRHQX1 reg_in_plain_key_out_reg_26_ ( .D(reg_in_n286), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[26]) );
  DFFRHQX1 reg_in_plain_key_out_reg_27_ ( .D(reg_in_n287), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[27]) );
  DFFRHQX1 reg_in_plain_key_out_reg_28_ ( .D(reg_in_n288), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[28]) );
  DFFRHQX1 reg_in_plain_key_out_reg_29_ ( .D(reg_in_n289), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[29]) );
  DFFRHQX1 reg_in_plain_key_out_reg_30_ ( .D(reg_in_n290), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[30]) );
  DFFRHQX1 reg_in_plain_key_out_reg_31_ ( .D(reg_in_n291), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[31]) );
  DFFRHQX1 reg_in_plain_key_out_reg_56_ ( .D(reg_in_n316), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[56]) );
  DFFRHQX1 reg_in_plain_key_out_reg_57_ ( .D(reg_in_n317), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[57]) );
  DFFRHQX1 reg_in_plain_key_out_reg_58_ ( .D(reg_in_n318), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[58]) );
  DFFRHQX1 reg_in_plain_key_out_reg_59_ ( .D(reg_in_n319), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[59]) );
  DFFRHQX1 reg_in_plain_key_out_reg_60_ ( .D(reg_in_n320), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[60]) );
  DFFRHQX1 reg_in_plain_key_out_reg_61_ ( .D(reg_in_n321), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[61]) );
  DFFRHQX1 reg_in_plain_key_out_reg_62_ ( .D(reg_in_n322), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[62]) );
  DFFRHQX1 reg_in_plain_key_out_reg_63_ ( .D(reg_in_n323), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[63]) );
  DFFRHQX1 reg_in_plain_key_out_reg_88_ ( .D(reg_in_n348), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[88]) );
  DFFRHQX1 reg_in_plain_key_out_reg_89_ ( .D(reg_in_n349), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[89]) );
  DFFRHQX1 reg_in_plain_key_out_reg_90_ ( .D(reg_in_n350), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[90]) );
  DFFRHQX1 reg_in_plain_key_out_reg_91_ ( .D(reg_in_n351), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[91]) );
  DFFRHQX1 reg_in_plain_key_out_reg_92_ ( .D(reg_in_n352), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[92]) );
  DFFRHQX1 reg_in_plain_key_out_reg_93_ ( .D(reg_in_n353), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[93]) );
  DFFRHQX1 reg_in_plain_key_out_reg_94_ ( .D(reg_in_n354), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[94]) );
  DFFRHQX1 reg_in_plain_key_out_reg_95_ ( .D(reg_in_n355), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[95]) );
  DFFRHQX1 reg_in_plain_key_out_reg_120_ ( .D(reg_in_n380), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[120]) );
  DFFRHQX1 reg_in_plain_key_out_reg_121_ ( .D(reg_in_n381), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[121]) );
  DFFRHQX1 reg_in_plain_key_out_reg_122_ ( .D(reg_in_n382), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[122]) );
  DFFRHQX1 reg_in_plain_key_out_reg_123_ ( .D(reg_in_n383), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[123]) );
  DFFRHQX1 reg_in_plain_key_out_reg_124_ ( .D(reg_in_n384), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[124]) );
  DFFRHQX1 reg_in_plain_key_out_reg_125_ ( .D(reg_in_n385), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[125]) );
  DFFRHQX1 reg_in_plain_key_out_reg_126_ ( .D(reg_in_n386), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[126]) );
  DFFRHQX1 reg_in_plain_key_out_reg_127_ ( .D(reg_in_n387), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[127]) );
  DFFRHQX1 reg_in_plain_key_out_reg_0_ ( .D(reg_in_n260), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[0]) );
  DFFRHQX1 reg_in_plain_key_out_reg_1_ ( .D(reg_in_n261), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[1]) );
  DFFRHQX1 reg_in_plain_key_out_reg_2_ ( .D(reg_in_n262), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[2]) );
  DFFRHQX1 reg_in_plain_key_out_reg_3_ ( .D(reg_in_n263), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[3]) );
  DFFRHQX1 reg_in_plain_key_out_reg_4_ ( .D(reg_in_n264), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[4]) );
  DFFRHQX1 reg_in_plain_key_out_reg_8_ ( .D(reg_in_n268), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[8]) );
  DFFRHQX1 reg_in_plain_key_out_reg_9_ ( .D(reg_in_n269), .CK(clk_48Mhz), .RN(
        reset_n), .Q(Din[9]) );
  DFFRHQX1 reg_in_plain_key_out_reg_10_ ( .D(reg_in_n270), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[10]) );
  DFFRHQX1 reg_in_plain_key_out_reg_11_ ( .D(reg_in_n271), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[11]) );
  DFFRHQX1 reg_in_plain_key_out_reg_12_ ( .D(reg_in_n272), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[12]) );
  DFFRHQX1 reg_in_plain_key_out_reg_13_ ( .D(reg_in_n273), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[13]) );
  DFFRHQX1 reg_in_plain_key_out_reg_14_ ( .D(reg_in_n274), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[14]) );
  DFFRHQX1 reg_in_plain_key_out_reg_15_ ( .D(reg_in_n275), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[15]) );
  DFFRHQX1 reg_in_plain_key_out_reg_16_ ( .D(reg_in_n276), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[16]) );
  DFFRHQX1 reg_in_plain_key_out_reg_17_ ( .D(reg_in_n277), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[17]) );
  DFFRHQX1 reg_in_plain_key_out_reg_18_ ( .D(reg_in_n278), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[18]) );
  DFFRHQX1 reg_in_plain_key_out_reg_19_ ( .D(reg_in_n279), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[19]) );
  DFFRHQX1 reg_in_plain_key_out_reg_20_ ( .D(reg_in_n280), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[20]) );
  DFFRHQX1 reg_in_plain_key_out_reg_21_ ( .D(reg_in_n281), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[21]) );
  DFFRHQX1 reg_in_plain_key_out_reg_22_ ( .D(reg_in_n282), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[22]) );
  DFFRHQX1 reg_in_plain_key_out_reg_23_ ( .D(reg_in_n283), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[23]) );
  DFFRHQX1 reg_in_plain_key_out_reg_32_ ( .D(reg_in_n292), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[32]) );
  DFFRHQX1 reg_in_plain_key_out_reg_33_ ( .D(reg_in_n293), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[33]) );
  DFFRHQX1 reg_in_plain_key_out_reg_34_ ( .D(reg_in_n294), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[34]) );
  DFFRHQX1 reg_in_plain_key_out_reg_35_ ( .D(reg_in_n295), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[35]) );
  DFFRHQX1 reg_in_plain_key_out_reg_36_ ( .D(reg_in_n296), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[36]) );
  DFFRHQX1 reg_in_plain_key_out_reg_37_ ( .D(reg_in_n297), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[37]) );
  DFFRHQX1 reg_in_plain_key_out_reg_38_ ( .D(reg_in_n298), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[38]) );
  DFFRHQX1 reg_in_plain_key_out_reg_39_ ( .D(reg_in_n299), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[39]) );
  DFFRHQX1 reg_in_plain_key_out_reg_40_ ( .D(reg_in_n300), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[40]) );
  DFFRHQX1 reg_in_plain_key_out_reg_41_ ( .D(reg_in_n301), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[41]) );
  DFFRHQX1 reg_in_plain_key_out_reg_42_ ( .D(reg_in_n302), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[42]) );
  DFFRHQX1 reg_in_plain_key_out_reg_43_ ( .D(reg_in_n303), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[43]) );
  DFFRHQX1 reg_in_plain_key_out_reg_44_ ( .D(reg_in_n304), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[44]) );
  DFFRHQX1 reg_in_plain_key_out_reg_45_ ( .D(reg_in_n305), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[45]) );
  DFFRHQX1 reg_in_plain_key_out_reg_46_ ( .D(reg_in_n306), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[46]) );
  DFFRHQX1 reg_in_plain_key_out_reg_47_ ( .D(reg_in_n307), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[47]) );
  DFFRHQX1 reg_in_plain_key_out_reg_48_ ( .D(reg_in_n308), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[48]) );
  DFFRHQX1 reg_in_plain_key_out_reg_49_ ( .D(reg_in_n309), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[49]) );
  DFFRHQX1 reg_in_plain_key_out_reg_50_ ( .D(reg_in_n310), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[50]) );
  DFFRHQX1 reg_in_plain_key_out_reg_51_ ( .D(reg_in_n311), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[51]) );
  DFFRHQX1 reg_in_plain_key_out_reg_52_ ( .D(reg_in_n312), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[52]) );
  DFFRHQX1 reg_in_plain_key_out_reg_53_ ( .D(reg_in_n313), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[53]) );
  DFFRHQX1 reg_in_plain_key_out_reg_54_ ( .D(reg_in_n314), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[54]) );
  DFFRHQX1 reg_in_plain_key_out_reg_55_ ( .D(reg_in_n315), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[55]) );
  DFFRHQX1 reg_in_plain_key_out_reg_64_ ( .D(reg_in_n324), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[64]) );
  DFFRHQX1 reg_in_plain_key_out_reg_65_ ( .D(reg_in_n325), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[65]) );
  DFFRHQX1 reg_in_plain_key_out_reg_66_ ( .D(reg_in_n326), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[66]) );
  DFFRHQX1 reg_in_plain_key_out_reg_67_ ( .D(reg_in_n327), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[67]) );
  DFFRHQX1 reg_in_plain_key_out_reg_68_ ( .D(reg_in_n328), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[68]) );
  DFFRHQX1 reg_in_plain_key_out_reg_69_ ( .D(reg_in_n329), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[69]) );
  DFFRHQX1 reg_in_plain_key_out_reg_70_ ( .D(reg_in_n330), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[70]) );
  DFFRHQX1 reg_in_plain_key_out_reg_71_ ( .D(reg_in_n331), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[71]) );
  DFFRHQX1 reg_in_plain_key_out_reg_72_ ( .D(reg_in_n332), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[72]) );
  DFFRHQX1 reg_in_plain_key_out_reg_73_ ( .D(reg_in_n333), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[73]) );
  DFFRHQX1 reg_in_plain_key_out_reg_74_ ( .D(reg_in_n334), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[74]) );
  DFFRHQX1 reg_in_plain_key_out_reg_76_ ( .D(reg_in_n336), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[76]) );
  DFFRHQX1 reg_in_plain_key_out_reg_77_ ( .D(reg_in_n337), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[77]) );
  DFFRHQX1 reg_in_plain_key_out_reg_78_ ( .D(reg_in_n338), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[78]) );
  DFFRHQX1 reg_in_plain_key_out_reg_79_ ( .D(reg_in_n339), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[79]) );
  DFFRHQX1 reg_in_plain_key_out_reg_80_ ( .D(reg_in_n340), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[80]) );
  DFFRHQX1 reg_in_plain_key_out_reg_81_ ( .D(reg_in_n341), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[81]) );
  DFFRHQX1 reg_in_plain_key_out_reg_82_ ( .D(reg_in_n342), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[82]) );
  DFFRHQX1 reg_in_plain_key_out_reg_83_ ( .D(reg_in_n343), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[83]) );
  DFFRHQX1 reg_in_plain_key_out_reg_84_ ( .D(reg_in_n344), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[84]) );
  DFFRHQX1 reg_in_plain_key_out_reg_85_ ( .D(reg_in_n345), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[85]) );
  DFFRHQX1 reg_in_plain_key_out_reg_86_ ( .D(reg_in_n346), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[86]) );
  DFFRHQX1 reg_in_plain_key_out_reg_87_ ( .D(reg_in_n347), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[87]) );
  DFFRHQX1 reg_in_plain_key_out_reg_96_ ( .D(reg_in_n356), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[96]) );
  DFFRHQX1 reg_in_plain_key_out_reg_97_ ( .D(reg_in_n357), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[97]) );
  DFFRHQX1 reg_in_plain_key_out_reg_98_ ( .D(reg_in_n358), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[98]) );
  DFFRHQX1 reg_in_plain_key_out_reg_99_ ( .D(reg_in_n359), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[99]) );
  DFFRHQX1 reg_in_plain_key_out_reg_100_ ( .D(reg_in_n360), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[100]) );
  DFFRHQX1 reg_in_plain_key_out_reg_101_ ( .D(reg_in_n361), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[101]) );
  DFFRHQX1 reg_in_plain_key_out_reg_102_ ( .D(reg_in_n362), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[102]) );
  DFFRHQX1 reg_in_plain_key_out_reg_103_ ( .D(reg_in_n363), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[103]) );
  DFFRHQX1 reg_in_plain_key_out_reg_104_ ( .D(reg_in_n364), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[104]) );
  DFFRHQX1 reg_in_plain_key_out_reg_105_ ( .D(reg_in_n365), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[105]) );
  DFFRHQX1 reg_in_plain_key_out_reg_106_ ( .D(reg_in_n366), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[106]) );
  DFFRHQX1 reg_in_plain_key_out_reg_107_ ( .D(reg_in_n367), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[107]) );
  DFFRHQX1 reg_in_plain_key_out_reg_108_ ( .D(reg_in_n368), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[108]) );
  DFFRHQX1 reg_in_plain_key_out_reg_109_ ( .D(reg_in_n369), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[109]) );
  DFFRHQX1 reg_in_plain_key_out_reg_110_ ( .D(reg_in_n370), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[110]) );
  DFFRHQX1 reg_in_plain_key_out_reg_111_ ( .D(reg_in_n371), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[111]) );
  DFFRHQX1 reg_in_plain_key_out_reg_112_ ( .D(reg_in_n372), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[112]) );
  DFFRHQX1 reg_in_plain_key_out_reg_113_ ( .D(reg_in_n373), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[113]) );
  DFFRHQX1 reg_in_plain_key_out_reg_114_ ( .D(reg_in_n374), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[114]) );
  DFFRHQX1 reg_in_plain_key_out_reg_115_ ( .D(reg_in_n375), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[115]) );
  DFFRHQX1 reg_in_plain_key_out_reg_116_ ( .D(reg_in_n376), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[116]) );
  DFFRHQX1 reg_in_plain_key_out_reg_117_ ( .D(reg_in_n377), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[117]) );
  DFFRHQX1 reg_in_plain_key_out_reg_118_ ( .D(reg_in_n378), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[118]) );
  DFFRHQX1 reg_in_plain_key_out_reg_119_ ( .D(reg_in_n379), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[119]) );
  DFFRHQX1 reg_in_plain_key_out_reg_128_ ( .D(reg_in_n388), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[128]) );
  DFFRHQX1 reg_in_plain_key_out_reg_129_ ( .D(reg_in_n389), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[129]) );
  DFFRHQX1 reg_in_plain_key_out_reg_130_ ( .D(reg_in_n390), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[130]) );
  DFFRHQX1 reg_in_plain_key_out_reg_131_ ( .D(reg_in_n391), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[131]) );
  DFFRHQX1 reg_in_plain_key_out_reg_132_ ( .D(reg_in_n392), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[132]) );
  DFFRHQX1 reg_in_plain_key_out_reg_133_ ( .D(reg_in_n393), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[133]) );
  DFFRHQX1 reg_in_plain_key_out_reg_134_ ( .D(reg_in_n394), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[134]) );
  DFFRHQX1 reg_in_plain_key_out_reg_135_ ( .D(reg_in_n395), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[135]) );
  DFFRHQX1 reg_in_plain_key_out_reg_136_ ( .D(reg_in_n396), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[136]) );
  DFFRHQX1 reg_in_plain_key_out_reg_137_ ( .D(reg_in_n397), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[137]) );
  DFFRHQX1 reg_in_plain_key_out_reg_138_ ( .D(reg_in_n398), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[138]) );
  DFFRHQX1 reg_in_plain_key_out_reg_139_ ( .D(reg_in_n399), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[139]) );
  DFFRHQX1 reg_in_plain_key_out_reg_140_ ( .D(reg_in_n400), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[140]) );
  DFFRHQX1 reg_in_plain_key_out_reg_141_ ( .D(reg_in_n401), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[141]) );
  DFFRHQX1 reg_in_plain_key_out_reg_142_ ( .D(reg_in_n402), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[142]) );
  DFFRHQX1 reg_in_plain_key_out_reg_143_ ( .D(reg_in_n403), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[143]) );
  DFFRHQX1 reg_in_plain_key_out_reg_144_ ( .D(reg_in_n404), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[144]) );
  DFFRHQX1 reg_in_plain_key_out_reg_145_ ( .D(reg_in_n405), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[145]) );
  DFFRHQX1 reg_in_plain_key_out_reg_146_ ( .D(reg_in_n406), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[146]) );
  DFFRHQX1 reg_in_plain_key_out_reg_147_ ( .D(reg_in_n407), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[147]) );
  DFFRHQX1 reg_in_plain_key_out_reg_148_ ( .D(reg_in_n408), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[148]) );
  DFFRHQX1 reg_in_plain_key_out_reg_149_ ( .D(reg_in_n409), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[149]) );
  DFFRHQX1 reg_in_plain_key_out_reg_150_ ( .D(reg_in_n410), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[150]) );
  DFFRHQX1 reg_in_plain_key_out_reg_151_ ( .D(reg_in_n411), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[151]) );
  DFFRHQX1 reg_in_plain_key_out_reg_152_ ( .D(reg_in_n412), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[152]) );
  DFFRHQX1 reg_in_plain_key_out_reg_153_ ( .D(reg_in_n413), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[153]) );
  DFFRHQX1 reg_in_plain_key_out_reg_154_ ( .D(reg_in_n414), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[154]) );
  DFFRHQX1 reg_in_plain_key_out_reg_155_ ( .D(reg_in_n415), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[155]) );
  DFFRHQX1 reg_in_plain_key_out_reg_156_ ( .D(reg_in_n416), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[156]) );
  DFFRHQX1 reg_in_plain_key_out_reg_157_ ( .D(reg_in_n417), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[157]) );
  DFFRHQX1 reg_in_plain_key_out_reg_158_ ( .D(reg_in_n418), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[158]) );
  DFFRHQX1 reg_in_plain_key_out_reg_159_ ( .D(reg_in_n419), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[159]) );
  DFFRHQX1 reg_in_plain_key_out_reg_160_ ( .D(reg_in_n420), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[160]) );
  DFFRHQX1 reg_in_plain_key_out_reg_161_ ( .D(reg_in_n421), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[161]) );
  DFFRHQX1 reg_in_plain_key_out_reg_162_ ( .D(reg_in_n422), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[162]) );
  DFFRHQX1 reg_in_plain_key_out_reg_163_ ( .D(reg_in_n423), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[163]) );
  DFFRHQX1 reg_in_plain_key_out_reg_164_ ( .D(reg_in_n424), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[164]) );
  DFFRHQX1 reg_in_plain_key_out_reg_165_ ( .D(reg_in_n425), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[165]) );
  DFFRHQX1 reg_in_plain_key_out_reg_166_ ( .D(reg_in_n426), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[166]) );
  DFFRHQX1 reg_in_plain_key_out_reg_167_ ( .D(reg_in_n427), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[167]) );
  DFFRHQX1 reg_in_plain_key_out_reg_168_ ( .D(reg_in_n428), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[168]) );
  DFFRHQX1 reg_in_plain_key_out_reg_169_ ( .D(reg_in_n429), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[169]) );
  DFFRHQX1 reg_in_plain_key_out_reg_170_ ( .D(reg_in_n430), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[170]) );
  DFFRHQX1 reg_in_plain_key_out_reg_171_ ( .D(reg_in_n431), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[171]) );
  DFFRHQX1 reg_in_plain_key_out_reg_172_ ( .D(reg_in_n432), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[172]) );
  DFFRHQX1 reg_in_plain_key_out_reg_173_ ( .D(reg_in_n433), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[173]) );
  DFFRHQX1 reg_in_plain_key_out_reg_174_ ( .D(reg_in_n434), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[174]) );
  DFFRHQX1 reg_in_plain_key_out_reg_175_ ( .D(reg_in_n435), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[175]) );
  DFFRHQX1 reg_in_plain_key_out_reg_176_ ( .D(reg_in_n436), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[176]) );
  DFFRHQX1 reg_in_plain_key_out_reg_177_ ( .D(reg_in_n437), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[177]) );
  DFFRHQX1 reg_in_plain_key_out_reg_178_ ( .D(reg_in_n438), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[178]) );
  DFFRHQX1 reg_in_plain_key_out_reg_179_ ( .D(reg_in_n439), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[179]) );
  DFFRHQX1 reg_in_plain_key_out_reg_180_ ( .D(reg_in_n440), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[180]) );
  DFFRHQX1 reg_in_plain_key_out_reg_181_ ( .D(reg_in_n441), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[181]) );
  DFFRHQX1 reg_in_plain_key_out_reg_182_ ( .D(reg_in_n442), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[182]) );
  DFFRHQX1 reg_in_plain_key_out_reg_183_ ( .D(reg_in_n443), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[183]) );
  DFFRHQX1 reg_in_plain_key_out_reg_184_ ( .D(reg_in_n444), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[184]) );
  DFFRHQX1 reg_in_plain_key_out_reg_185_ ( .D(reg_in_n445), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[185]) );
  DFFRHQX1 reg_in_plain_key_out_reg_186_ ( .D(reg_in_n446), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[186]) );
  DFFRHQX1 reg_in_plain_key_out_reg_187_ ( .D(reg_in_n447), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[187]) );
  DFFRHQX1 reg_in_plain_key_out_reg_188_ ( .D(reg_in_n448), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[188]) );
  DFFRHQX1 reg_in_plain_key_out_reg_189_ ( .D(reg_in_n449), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[189]) );
  DFFRHQX1 reg_in_plain_key_out_reg_190_ ( .D(reg_in_n450), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[190]) );
  DFFRHQX1 reg_in_plain_key_out_reg_191_ ( .D(reg_in_n451), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[191]) );
  DFFRHQX1 reg_in_plain_key_out_reg_192_ ( .D(reg_in_n452), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[192]) );
  DFFRHQX1 reg_in_plain_key_out_reg_193_ ( .D(reg_in_n453), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[193]) );
  DFFRHQX1 reg_in_plain_key_out_reg_194_ ( .D(reg_in_n454), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[194]) );
  DFFRHQX1 reg_in_plain_key_out_reg_195_ ( .D(reg_in_n455), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[195]) );
  DFFRHQX1 reg_in_plain_key_out_reg_196_ ( .D(reg_in_n456), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[196]) );
  DFFRHQX1 reg_in_plain_key_out_reg_197_ ( .D(reg_in_n457), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[197]) );
  DFFRHQX1 reg_in_plain_key_out_reg_198_ ( .D(reg_in_n458), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[198]) );
  DFFRHQX1 reg_in_plain_key_out_reg_199_ ( .D(reg_in_n459), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[199]) );
  DFFRHQX1 reg_in_plain_key_out_reg_200_ ( .D(reg_in_n460), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[200]) );
  DFFRHQX1 reg_in_plain_key_out_reg_201_ ( .D(reg_in_n461), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[201]) );
  DFFRHQX1 reg_in_plain_key_out_reg_202_ ( .D(reg_in_n462), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[202]) );
  DFFRHQX1 reg_in_plain_key_out_reg_203_ ( .D(reg_in_n463), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[203]) );
  DFFRHQX1 reg_in_plain_key_out_reg_204_ ( .D(reg_in_n464), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[204]) );
  DFFRHQX1 reg_in_plain_key_out_reg_205_ ( .D(reg_in_n465), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[205]) );
  DFFRHQX1 reg_in_plain_key_out_reg_206_ ( .D(reg_in_n466), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[206]) );
  DFFRHQX1 reg_in_plain_key_out_reg_207_ ( .D(reg_in_n467), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[207]) );
  DFFRHQX1 reg_in_plain_key_out_reg_208_ ( .D(reg_in_n468), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[208]) );
  DFFRHQX1 reg_in_plain_key_out_reg_209_ ( .D(reg_in_n469), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[209]) );
  DFFRHQX1 reg_in_plain_key_out_reg_210_ ( .D(reg_in_n470), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[210]) );
  DFFRHQX1 reg_in_plain_key_out_reg_211_ ( .D(reg_in_n471), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[211]) );
  DFFRHQX1 reg_in_plain_key_out_reg_212_ ( .D(reg_in_n472), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[212]) );
  DFFRHQX1 reg_in_plain_key_out_reg_213_ ( .D(reg_in_n473), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[213]) );
  DFFRHQX1 reg_in_plain_key_out_reg_214_ ( .D(reg_in_n474), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[214]) );
  DFFRHQX1 reg_in_plain_key_out_reg_215_ ( .D(reg_in_n475), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[215]) );
  DFFRHQX1 reg_in_plain_key_out_reg_216_ ( .D(reg_in_n476), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[216]) );
  DFFRHQX1 reg_in_plain_key_out_reg_217_ ( .D(reg_in_n477), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[217]) );
  DFFRHQX1 reg_in_plain_key_out_reg_218_ ( .D(reg_in_n478), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(Din[218]) );
  DFFRHQX1 reg_in_plain_text_reg_240_ ( .D(reg_in_n517), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[240]) );
  DFFRHQX1 reg_in_plain_text_reg_232_ ( .D(reg_in_n518), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[232]) );
  DFFRHQX1 reg_in_plain_text_reg_224_ ( .D(reg_in_n519), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[224]) );
  DFFRHQX1 reg_in_plain_text_reg_216_ ( .D(reg_in_n520), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[216]) );
  DFFRHQX1 reg_in_plain_text_reg_208_ ( .D(reg_in_n521), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[208]) );
  DFFRHQX1 reg_in_plain_text_reg_200_ ( .D(reg_in_n522), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[200]) );
  DFFRHQX1 reg_in_plain_text_reg_192_ ( .D(reg_in_n523), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[192]) );
  DFFRHQX1 reg_in_plain_text_reg_184_ ( .D(reg_in_n524), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[184]) );
  DFFRHQX1 reg_in_plain_text_reg_176_ ( .D(reg_in_n525), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[176]) );
  DFFRHQX1 reg_in_plain_text_reg_168_ ( .D(reg_in_n526), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[168]) );
  DFFRHQX1 reg_in_plain_text_reg_160_ ( .D(reg_in_n527), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[160]) );
  DFFRHQX1 reg_in_plain_text_reg_152_ ( .D(reg_in_n528), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[152]) );
  DFFRHQX1 reg_in_plain_text_reg_144_ ( .D(reg_in_n529), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[144]) );
  DFFRHQX1 reg_in_plain_text_reg_136_ ( .D(reg_in_n530), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[136]) );
  DFFRHQX1 reg_in_plain_text_reg_128_ ( .D(reg_in_n531), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[128]) );
  DFFRHQX1 reg_in_plain_text_reg_120_ ( .D(reg_in_n532), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[120]) );
  DFFRHQX1 reg_in_plain_text_reg_112_ ( .D(reg_in_n533), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[112]) );
  DFFRHQX1 reg_in_plain_text_reg_104_ ( .D(reg_in_n534), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[104]) );
  DFFRHQX1 reg_in_plain_text_reg_96_ ( .D(reg_in_n535), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[96]) );
  DFFRHQX1 reg_in_plain_text_reg_88_ ( .D(reg_in_n536), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[88]) );
  DFFRHQX1 reg_in_plain_text_reg_80_ ( .D(reg_in_n537), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[80]) );
  DFFRHQX1 reg_in_plain_text_reg_72_ ( .D(reg_in_n538), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[72]) );
  DFFRHQX1 reg_in_plain_text_reg_64_ ( .D(reg_in_n539), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[64]) );
  DFFRHQX1 reg_in_plain_text_reg_56_ ( .D(reg_in_n540), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[56]) );
  DFFRHQX1 reg_in_plain_text_reg_48_ ( .D(reg_in_n541), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[48]) );
  DFFRHQX1 reg_in_plain_text_reg_40_ ( .D(reg_in_n542), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[40]) );
  DFFRHQX1 reg_in_plain_text_reg_32_ ( .D(reg_in_n543), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[32]) );
  DFFRHQX1 reg_in_plain_text_reg_24_ ( .D(reg_in_n544), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[24]) );
  DFFRHQX1 reg_in_plain_text_reg_16_ ( .D(reg_in_n545), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[16]) );
  DFFRHQX1 reg_in_plain_text_reg_8_ ( .D(reg_in_n546), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[8]) );
  DFFRHQX1 reg_in_plain_text_reg_0_ ( .D(reg_in_n547), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[0]) );
  DFFRHQX1 reg_in_plain_text_reg_241_ ( .D(reg_in_n549), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[241]) );
  DFFRHQX1 reg_in_plain_text_reg_233_ ( .D(reg_in_n550), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[233]) );
  DFFRHQX1 reg_in_plain_text_reg_225_ ( .D(reg_in_n551), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[225]) );
  DFFRHQX1 reg_in_plain_text_reg_217_ ( .D(reg_in_n552), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[217]) );
  DFFRHQX1 reg_in_plain_text_reg_209_ ( .D(reg_in_n553), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[209]) );
  DFFRHQX1 reg_in_plain_text_reg_201_ ( .D(reg_in_n554), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[201]) );
  DFFRHQX1 reg_in_plain_text_reg_193_ ( .D(reg_in_n555), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[193]) );
  DFFRHQX1 reg_in_plain_text_reg_185_ ( .D(reg_in_n556), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[185]) );
  DFFRHQX1 reg_in_plain_text_reg_177_ ( .D(reg_in_n557), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[177]) );
  DFFRHQX1 reg_in_plain_text_reg_169_ ( .D(reg_in_n558), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[169]) );
  DFFRHQX1 reg_in_plain_text_reg_161_ ( .D(reg_in_n559), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[161]) );
  DFFRHQX1 reg_in_plain_text_reg_153_ ( .D(reg_in_n560), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[153]) );
  DFFRHQX1 reg_in_plain_text_reg_145_ ( .D(reg_in_n561), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[145]) );
  DFFRHQX1 reg_in_plain_text_reg_137_ ( .D(reg_in_n562), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[137]) );
  DFFRHQX1 reg_in_plain_text_reg_129_ ( .D(reg_in_n563), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[129]) );
  DFFRHQX1 reg_in_plain_text_reg_121_ ( .D(reg_in_n564), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[121]) );
  DFFRHQX1 reg_in_plain_text_reg_113_ ( .D(reg_in_n565), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[113]) );
  DFFRHQX1 reg_in_plain_text_reg_105_ ( .D(reg_in_n566), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[105]) );
  DFFRHQX1 reg_in_plain_text_reg_97_ ( .D(reg_in_n567), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[97]) );
  DFFRHQX1 reg_in_plain_text_reg_89_ ( .D(reg_in_n568), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[89]) );
  DFFRHQX1 reg_in_plain_text_reg_81_ ( .D(reg_in_n569), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[81]) );
  DFFRHQX1 reg_in_plain_text_reg_73_ ( .D(reg_in_n570), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[73]) );
  DFFRHQX1 reg_in_plain_text_reg_65_ ( .D(reg_in_n571), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[65]) );
  DFFRHQX1 reg_in_plain_text_reg_57_ ( .D(reg_in_n572), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[57]) );
  DFFRHQX1 reg_in_plain_text_reg_49_ ( .D(reg_in_n573), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[49]) );
  DFFRHQX1 reg_in_plain_text_reg_41_ ( .D(reg_in_n574), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[41]) );
  DFFRHQX1 reg_in_plain_text_reg_33_ ( .D(reg_in_n575), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[33]) );
  DFFRHQX1 reg_in_plain_text_reg_25_ ( .D(reg_in_n576), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[25]) );
  DFFRHQX1 reg_in_plain_text_reg_17_ ( .D(reg_in_n577), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[17]) );
  DFFRHQX1 reg_in_plain_text_reg_9_ ( .D(reg_in_n578), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[9]) );
  DFFRHQX1 reg_in_plain_text_reg_1_ ( .D(reg_in_n579), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[1]) );
  DFFRHQX1 reg_in_plain_text_reg_242_ ( .D(reg_in_n581), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[242]) );
  DFFRHQX1 reg_in_plain_text_reg_234_ ( .D(reg_in_n582), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[234]) );
  DFFRHQX1 reg_in_plain_text_reg_226_ ( .D(reg_in_n583), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[226]) );
  DFFRHQX1 reg_in_plain_text_reg_218_ ( .D(reg_in_n584), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[218]) );
  DFFRHQX1 reg_in_plain_text_reg_210_ ( .D(reg_in_n585), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[210]) );
  DFFRHQX1 reg_in_plain_text_reg_202_ ( .D(reg_in_n586), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[202]) );
  DFFRHQX1 reg_in_plain_text_reg_194_ ( .D(reg_in_n587), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[194]) );
  DFFRHQX1 reg_in_plain_text_reg_186_ ( .D(reg_in_n588), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[186]) );
  DFFRHQX1 reg_in_plain_text_reg_178_ ( .D(reg_in_n589), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[178]) );
  DFFRHQX1 reg_in_plain_text_reg_170_ ( .D(reg_in_n590), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[170]) );
  DFFRHQX1 reg_in_plain_text_reg_162_ ( .D(reg_in_n591), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[162]) );
  DFFRHQX1 reg_in_plain_text_reg_154_ ( .D(reg_in_n592), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[154]) );
  DFFRHQX1 reg_in_plain_text_reg_146_ ( .D(reg_in_n593), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[146]) );
  DFFRHQX1 reg_in_plain_text_reg_138_ ( .D(reg_in_n594), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[138]) );
  DFFRHQX1 reg_in_plain_text_reg_130_ ( .D(reg_in_n595), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[130]) );
  DFFRHQX1 reg_in_plain_text_reg_122_ ( .D(reg_in_n596), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[122]) );
  DFFRHQX1 reg_in_plain_text_reg_114_ ( .D(reg_in_n597), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[114]) );
  DFFRHQX1 reg_in_plain_text_reg_106_ ( .D(reg_in_n598), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[106]) );
  DFFRHQX1 reg_in_plain_text_reg_98_ ( .D(reg_in_n599), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[98]) );
  DFFRHQX1 reg_in_plain_text_reg_90_ ( .D(reg_in_n600), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[90]) );
  DFFRHQX1 reg_in_plain_text_reg_82_ ( .D(reg_in_n601), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[82]) );
  DFFRHQX1 reg_in_plain_text_reg_74_ ( .D(reg_in_n602), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[74]) );
  DFFRHQX1 reg_in_plain_text_reg_66_ ( .D(reg_in_n603), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[66]) );
  DFFRHQX1 reg_in_plain_text_reg_58_ ( .D(reg_in_n604), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[58]) );
  DFFRHQX1 reg_in_plain_text_reg_50_ ( .D(reg_in_n605), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[50]) );
  DFFRHQX1 reg_in_plain_text_reg_42_ ( .D(reg_in_n606), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[42]) );
  DFFRHQX1 reg_in_plain_text_reg_34_ ( .D(reg_in_n607), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[34]) );
  DFFRHQX1 reg_in_plain_text_reg_26_ ( .D(reg_in_n608), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[26]) );
  DFFRHQX1 reg_in_plain_text_reg_18_ ( .D(reg_in_n609), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[18]) );
  DFFRHQX1 reg_in_plain_text_reg_10_ ( .D(reg_in_n610), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[10]) );
  DFFRHQX1 reg_in_plain_text_reg_2_ ( .D(reg_in_n611), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[2]) );
  DFFRHQX1 reg_in_plain_text_reg_243_ ( .D(reg_in_n613), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[243]) );
  DFFRHQX1 reg_in_plain_text_reg_235_ ( .D(reg_in_n614), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[235]) );
  DFFRHQX1 reg_in_plain_text_reg_227_ ( .D(reg_in_n615), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[227]) );
  DFFRHQX1 reg_in_plain_text_reg_219_ ( .D(reg_in_n616), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[219]) );
  DFFRHQX1 reg_in_plain_text_reg_211_ ( .D(reg_in_n617), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[211]) );
  DFFRHQX1 reg_in_plain_text_reg_203_ ( .D(reg_in_n618), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[203]) );
  DFFRHQX1 reg_in_plain_text_reg_195_ ( .D(reg_in_n619), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[195]) );
  DFFRHQX1 reg_in_plain_text_reg_187_ ( .D(reg_in_n620), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[187]) );
  DFFRHQX1 reg_in_plain_text_reg_179_ ( .D(reg_in_n621), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[179]) );
  DFFRHQX1 reg_in_plain_text_reg_171_ ( .D(reg_in_n622), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[171]) );
  DFFRHQX1 reg_in_plain_text_reg_163_ ( .D(reg_in_n623), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[163]) );
  DFFRHQX1 reg_in_plain_text_reg_155_ ( .D(reg_in_n624), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[155]) );
  DFFRHQX1 reg_in_plain_text_reg_147_ ( .D(reg_in_n625), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[147]) );
  DFFRHQX1 reg_in_plain_text_reg_139_ ( .D(reg_in_n626), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[139]) );
  DFFRHQX1 reg_in_plain_text_reg_131_ ( .D(reg_in_n627), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[131]) );
  DFFRHQX1 reg_in_plain_text_reg_123_ ( .D(reg_in_n628), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[123]) );
  DFFRHQX1 reg_in_plain_text_reg_115_ ( .D(reg_in_n629), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[115]) );
  DFFRHQX1 reg_in_plain_text_reg_107_ ( .D(reg_in_n630), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[107]) );
  DFFRHQX1 reg_in_plain_text_reg_99_ ( .D(reg_in_n631), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[99]) );
  DFFRHQX1 reg_in_plain_text_reg_91_ ( .D(reg_in_n632), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[91]) );
  DFFRHQX1 reg_in_plain_text_reg_83_ ( .D(reg_in_n633), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[83]) );
  DFFRHQX1 reg_in_plain_text_reg_75_ ( .D(reg_in_n634), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[75]) );
  DFFRHQX1 reg_in_plain_text_reg_67_ ( .D(reg_in_n635), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[67]) );
  DFFRHQX1 reg_in_plain_text_reg_59_ ( .D(reg_in_n636), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[59]) );
  DFFRHQX1 reg_in_plain_text_reg_51_ ( .D(reg_in_n637), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[51]) );
  DFFRHQX1 reg_in_plain_text_reg_43_ ( .D(reg_in_n638), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[43]) );
  DFFRHQX1 reg_in_plain_text_reg_35_ ( .D(reg_in_n639), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[35]) );
  DFFRHQX1 reg_in_plain_text_reg_27_ ( .D(reg_in_n640), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[27]) );
  DFFRHQX1 reg_in_plain_text_reg_19_ ( .D(reg_in_n641), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[19]) );
  DFFRHQX1 reg_in_plain_text_reg_11_ ( .D(reg_in_n642), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[11]) );
  DFFRHQX1 reg_in_plain_text_reg_3_ ( .D(reg_in_n643), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[3]) );
  DFFRHQX1 reg_in_plain_text_reg_244_ ( .D(reg_in_n645), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[244]) );
  DFFRHQX1 reg_in_plain_text_reg_236_ ( .D(reg_in_n646), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[236]) );
  DFFRHQX1 reg_in_plain_text_reg_228_ ( .D(reg_in_n647), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[228]) );
  DFFRHQX1 reg_in_plain_text_reg_220_ ( .D(reg_in_n648), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[220]) );
  DFFRHQX1 reg_in_plain_text_reg_212_ ( .D(reg_in_n649), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[212]) );
  DFFRHQX1 reg_in_plain_text_reg_204_ ( .D(reg_in_n650), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[204]) );
  DFFRHQX1 reg_in_plain_text_reg_196_ ( .D(reg_in_n651), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[196]) );
  DFFRHQX1 reg_in_plain_text_reg_188_ ( .D(reg_in_n652), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[188]) );
  DFFRHQX1 reg_in_plain_text_reg_180_ ( .D(reg_in_n653), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[180]) );
  DFFRHQX1 reg_in_plain_text_reg_172_ ( .D(reg_in_n654), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[172]) );
  DFFRHQX1 reg_in_plain_text_reg_164_ ( .D(reg_in_n655), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[164]) );
  DFFRHQX1 reg_in_plain_text_reg_156_ ( .D(reg_in_n656), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[156]) );
  DFFRHQX1 reg_in_plain_text_reg_148_ ( .D(reg_in_n657), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[148]) );
  DFFRHQX1 reg_in_plain_text_reg_140_ ( .D(reg_in_n658), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[140]) );
  DFFRHQX1 reg_in_plain_text_reg_132_ ( .D(reg_in_n659), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[132]) );
  DFFRHQX1 reg_in_plain_text_reg_124_ ( .D(reg_in_n660), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[124]) );
  DFFRHQX1 reg_in_plain_text_reg_116_ ( .D(reg_in_n661), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[116]) );
  DFFRHQX1 reg_in_plain_text_reg_108_ ( .D(reg_in_n662), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[108]) );
  DFFRHQX1 reg_in_plain_text_reg_100_ ( .D(reg_in_n663), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[100]) );
  DFFRHQX1 reg_in_plain_text_reg_92_ ( .D(reg_in_n664), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[92]) );
  DFFRHQX1 reg_in_plain_text_reg_84_ ( .D(reg_in_n665), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[84]) );
  DFFRHQX1 reg_in_plain_text_reg_76_ ( .D(reg_in_n666), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[76]) );
  DFFRHQX1 reg_in_plain_text_reg_68_ ( .D(reg_in_n667), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[68]) );
  DFFRHQX1 reg_in_plain_text_reg_60_ ( .D(reg_in_n668), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[60]) );
  DFFRHQX1 reg_in_plain_text_reg_52_ ( .D(reg_in_n669), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[52]) );
  DFFRHQX1 reg_in_plain_text_reg_44_ ( .D(reg_in_n670), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[44]) );
  DFFRHQX1 reg_in_plain_text_reg_36_ ( .D(reg_in_n671), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[36]) );
  DFFRHQX1 reg_in_plain_text_reg_28_ ( .D(reg_in_n672), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[28]) );
  DFFRHQX1 reg_in_plain_text_reg_20_ ( .D(reg_in_n673), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[20]) );
  DFFRHQX1 reg_in_plain_text_reg_12_ ( .D(reg_in_n674), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[12]) );
  DFFRHQX1 reg_in_plain_text_reg_4_ ( .D(reg_in_n675), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[4]) );
  DFFRHQX1 reg_in_plain_text_reg_245_ ( .D(reg_in_n677), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[245]) );
  DFFRHQX1 reg_in_plain_text_reg_237_ ( .D(reg_in_n678), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[237]) );
  DFFRHQX1 reg_in_plain_text_reg_229_ ( .D(reg_in_n679), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[229]) );
  DFFRHQX1 reg_in_plain_text_reg_221_ ( .D(reg_in_n680), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[221]) );
  DFFRHQX1 reg_in_plain_text_reg_213_ ( .D(reg_in_n681), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[213]) );
  DFFRHQX1 reg_in_plain_text_reg_205_ ( .D(reg_in_n682), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[205]) );
  DFFRHQX1 reg_in_plain_text_reg_197_ ( .D(reg_in_n683), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[197]) );
  DFFRHQX1 reg_in_plain_text_reg_189_ ( .D(reg_in_n684), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[189]) );
  DFFRHQX1 reg_in_plain_text_reg_181_ ( .D(reg_in_n685), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[181]) );
  DFFRHQX1 reg_in_plain_text_reg_173_ ( .D(reg_in_n686), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[173]) );
  DFFRHQX1 reg_in_plain_text_reg_165_ ( .D(reg_in_n687), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[165]) );
  DFFRHQX1 reg_in_plain_text_reg_157_ ( .D(reg_in_n688), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[157]) );
  DFFRHQX1 reg_in_plain_text_reg_149_ ( .D(reg_in_n689), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[149]) );
  DFFRHQX1 reg_in_plain_text_reg_141_ ( .D(reg_in_n690), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[141]) );
  DFFRHQX1 reg_in_plain_text_reg_133_ ( .D(reg_in_n691), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[133]) );
  DFFRHQX1 reg_in_plain_text_reg_125_ ( .D(reg_in_n692), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[125]) );
  DFFRHQX1 reg_in_plain_text_reg_117_ ( .D(reg_in_n693), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[117]) );
  DFFRHQX1 reg_in_plain_text_reg_109_ ( .D(reg_in_n694), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[109]) );
  DFFRHQX1 reg_in_plain_text_reg_101_ ( .D(reg_in_n695), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[101]) );
  DFFRHQX1 reg_in_plain_text_reg_93_ ( .D(reg_in_n696), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[93]) );
  DFFRHQX1 reg_in_plain_text_reg_85_ ( .D(reg_in_n697), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[85]) );
  DFFRHQX1 reg_in_plain_text_reg_77_ ( .D(reg_in_n698), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[77]) );
  DFFRHQX1 reg_in_plain_text_reg_69_ ( .D(reg_in_n699), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[69]) );
  DFFRHQX1 reg_in_plain_text_reg_61_ ( .D(reg_in_n700), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[61]) );
  DFFRHQX1 reg_in_plain_text_reg_53_ ( .D(reg_in_n701), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[53]) );
  DFFRHQX1 reg_in_plain_text_reg_45_ ( .D(reg_in_n702), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[45]) );
  DFFRHQX1 reg_in_plain_text_reg_37_ ( .D(reg_in_n703), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[37]) );
  DFFRHQX1 reg_in_plain_text_reg_29_ ( .D(reg_in_n704), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[29]) );
  DFFRHQX1 reg_in_plain_text_reg_21_ ( .D(reg_in_n705), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[21]) );
  DFFRHQX1 reg_in_plain_text_reg_13_ ( .D(reg_in_n706), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[13]) );
  DFFRHQX1 reg_in_plain_text_reg_5_ ( .D(reg_in_n707), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[5]) );
  DFFRHQX1 reg_in_plain_text_reg_246_ ( .D(reg_in_n709), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[246]) );
  DFFRHQX1 reg_in_plain_text_reg_238_ ( .D(reg_in_n710), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[238]) );
  DFFRHQX1 reg_in_plain_text_reg_230_ ( .D(reg_in_n711), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[230]) );
  DFFRHQX1 reg_in_plain_text_reg_222_ ( .D(reg_in_n712), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[222]) );
  DFFRHQX1 reg_in_plain_text_reg_214_ ( .D(reg_in_n713), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[214]) );
  DFFRHQX1 reg_in_plain_text_reg_206_ ( .D(reg_in_n714), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[206]) );
  DFFRHQX1 reg_in_plain_text_reg_198_ ( .D(reg_in_n715), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[198]) );
  DFFRHQX1 reg_in_plain_text_reg_190_ ( .D(reg_in_n716), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[190]) );
  DFFRHQX1 reg_in_plain_text_reg_182_ ( .D(reg_in_n717), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[182]) );
  DFFRHQX1 reg_in_plain_text_reg_174_ ( .D(reg_in_n718), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[174]) );
  DFFRHQX1 reg_in_plain_text_reg_166_ ( .D(reg_in_n719), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[166]) );
  DFFRHQX1 reg_in_plain_text_reg_158_ ( .D(reg_in_n720), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[158]) );
  DFFRHQX1 reg_in_plain_text_reg_150_ ( .D(reg_in_n721), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[150]) );
  DFFRHQX1 reg_in_plain_text_reg_142_ ( .D(reg_in_n722), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[142]) );
  DFFRHQX1 reg_in_plain_text_reg_134_ ( .D(reg_in_n723), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[134]) );
  DFFRHQX1 reg_in_plain_text_reg_126_ ( .D(reg_in_n724), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[126]) );
  DFFRHQX1 reg_in_plain_text_reg_118_ ( .D(reg_in_n725), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[118]) );
  DFFRHQX1 reg_in_plain_text_reg_110_ ( .D(reg_in_n726), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[110]) );
  DFFRHQX1 reg_in_plain_text_reg_102_ ( .D(reg_in_n727), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[102]) );
  DFFRHQX1 reg_in_plain_text_reg_94_ ( .D(reg_in_n728), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[94]) );
  DFFRHQX1 reg_in_plain_text_reg_86_ ( .D(reg_in_n729), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[86]) );
  DFFRHQX1 reg_in_plain_text_reg_78_ ( .D(reg_in_n730), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[78]) );
  DFFRHQX1 reg_in_plain_text_reg_70_ ( .D(reg_in_n731), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[70]) );
  DFFRHQX1 reg_in_plain_text_reg_62_ ( .D(reg_in_n732), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[62]) );
  DFFRHQX1 reg_in_plain_text_reg_54_ ( .D(reg_in_n733), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[54]) );
  DFFRHQX1 reg_in_plain_text_reg_46_ ( .D(reg_in_n734), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[46]) );
  DFFRHQX1 reg_in_plain_text_reg_38_ ( .D(reg_in_n735), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[38]) );
  DFFRHQX1 reg_in_plain_text_reg_30_ ( .D(reg_in_n736), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[30]) );
  DFFRHQX1 reg_in_plain_text_reg_22_ ( .D(reg_in_n737), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[22]) );
  DFFRHQX1 reg_in_plain_text_reg_14_ ( .D(reg_in_n738), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[14]) );
  DFFRHQX1 reg_in_plain_text_reg_6_ ( .D(reg_in_n739), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[6]) );
  DFFRHQX1 reg_in_plain_text_reg_247_ ( .D(reg_in_n741), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[247]) );
  DFFRHQX1 reg_in_plain_text_reg_239_ ( .D(reg_in_n742), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[239]) );
  DFFRHQX1 reg_in_plain_text_reg_231_ ( .D(reg_in_n743), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[231]) );
  DFFRHQX1 reg_in_plain_text_reg_223_ ( .D(reg_in_n744), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[223]) );
  DFFRHQX1 reg_in_plain_text_reg_215_ ( .D(reg_in_n745), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[215]) );
  DFFRHQX1 reg_in_plain_text_reg_207_ ( .D(reg_in_n746), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[207]) );
  DFFRHQX1 reg_in_plain_text_reg_199_ ( .D(reg_in_n747), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[199]) );
  DFFRHQX1 reg_in_plain_text_reg_191_ ( .D(reg_in_n748), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[191]) );
  DFFRHQX1 reg_in_plain_text_reg_183_ ( .D(reg_in_n749), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[183]) );
  DFFRHQX1 reg_in_plain_text_reg_175_ ( .D(reg_in_n750), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[175]) );
  DFFRHQX1 reg_in_plain_text_reg_167_ ( .D(reg_in_n751), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[167]) );
  DFFRHQX1 reg_in_plain_text_reg_159_ ( .D(reg_in_n752), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[159]) );
  DFFRHQX1 reg_in_plain_text_reg_151_ ( .D(reg_in_n753), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[151]) );
  DFFRHQX1 reg_in_plain_text_reg_143_ ( .D(reg_in_n754), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[143]) );
  DFFRHQX1 reg_in_plain_text_reg_135_ ( .D(reg_in_n755), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[135]) );
  DFFRHQX1 reg_in_plain_text_reg_127_ ( .D(reg_in_n756), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[127]) );
  DFFRHQX1 reg_in_plain_text_reg_119_ ( .D(reg_in_n757), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[119]) );
  DFFRHQX1 reg_in_plain_text_reg_111_ ( .D(reg_in_n758), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[111]) );
  DFFRHQX1 reg_in_plain_text_reg_103_ ( .D(reg_in_n759), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[103]) );
  DFFRHQX1 reg_in_plain_text_reg_95_ ( .D(reg_in_n760), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[95]) );
  DFFRHQX1 reg_in_plain_text_reg_87_ ( .D(reg_in_n761), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[87]) );
  DFFRHQX1 reg_in_plain_text_reg_79_ ( .D(reg_in_n762), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[79]) );
  DFFRHQX1 reg_in_plain_text_reg_71_ ( .D(reg_in_n763), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[71]) );
  DFFRHQX1 reg_in_plain_text_reg_63_ ( .D(reg_in_n764), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[63]) );
  DFFRHQX1 reg_in_plain_text_reg_55_ ( .D(reg_in_n765), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[55]) );
  DFFRHQX1 reg_in_plain_text_reg_47_ ( .D(reg_in_n766), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[47]) );
  DFFRHQX1 reg_in_plain_text_reg_39_ ( .D(reg_in_n767), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[39]) );
  DFFRHQX1 reg_in_plain_text_reg_31_ ( .D(reg_in_n768), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[31]) );
  DFFRHQX1 reg_in_plain_text_reg_23_ ( .D(reg_in_n769), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[23]) );
  DFFRHQX1 reg_in_plain_text_reg_15_ ( .D(reg_in_n770), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[15]) );
  DFFRHQX1 reg_in_plain_text_reg_7_ ( .D(reg_in_n771), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[7]) );
  DFFRHQX1 reg_in_plain_text_reg_248_ ( .D(reg_in_n516), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[248]) );
  DFFRHQX1 reg_in_plain_text_reg_249_ ( .D(reg_in_n548), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[249]) );
  DFFRHQX1 reg_in_plain_text_reg_250_ ( .D(reg_in_n580), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[250]) );
  DFFRHQX1 reg_in_plain_text_reg_251_ ( .D(reg_in_n612), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[251]) );
  DFFRHQX1 reg_in_plain_text_reg_252_ ( .D(reg_in_n644), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[252]) );
  DFFRHQX1 reg_in_plain_text_reg_253_ ( .D(reg_in_n676), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[253]) );
  DFFRHQX1 reg_in_plain_text_reg_254_ ( .D(reg_in_n708), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[254]) );
  DFFRHQX1 reg_in_plain_text_reg_255_ ( .D(reg_in_n740), .CK(clk_48Mhz), .RN(
        reset_n), .Q(reg_in_plain_text[255]) );
  INVX1 reg_out_U313 ( .A(reg_out_rdy0), .Y(reg_out_n310) );
  NOR2BX1 reg_out_U312 ( .AN(reg_out_rdy2), .B(reg_out_rdy1), .Y(
        cipher_byte_valid) );
  AOI22X1 reg_out_U311 ( .A0(reg_out_n280), .A1(reg_out_cipher_sample[126]), 
        .B0(cipher_byte_out[6]), .B1(reg_out_n2), .Y(reg_out_n16) );
  INVX1 reg_out_U310 ( .A(reg_out_n16), .Y(reg_out_n303) );
  AOI22X1 reg_out_U309 ( .A0(reg_out_n280), .A1(reg_out_cipher_sample[125]), 
        .B0(cipher_byte_out[5]), .B1(reg_out_n2), .Y(reg_out_n18) );
  INVX1 reg_out_U308 ( .A(reg_out_n18), .Y(reg_out_n304) );
  AOI22X1 reg_out_U307 ( .A0(reg_out_n280), .A1(reg_out_cipher_sample[124]), 
        .B0(cipher_byte_out[4]), .B1(reg_out_n2), .Y(reg_out_n20) );
  INVX1 reg_out_U306 ( .A(reg_out_n20), .Y(reg_out_n305) );
  AOI22X1 reg_out_U305 ( .A0(reg_out_n280), .A1(reg_out_cipher_sample[123]), 
        .B0(cipher_byte_out[3]), .B1(reg_out_n2), .Y(reg_out_n22) );
  INVX1 reg_out_U304 ( .A(reg_out_n22), .Y(reg_out_n306) );
  AOI22X1 reg_out_U303 ( .A0(reg_out_n3), .A1(reg_out_cipher_sample[122]), 
        .B0(cipher_byte_out[2]), .B1(reg_out_n2), .Y(reg_out_n24) );
  INVX1 reg_out_U302 ( .A(reg_out_n24), .Y(reg_out_n307) );
  AOI22X1 reg_out_U301 ( .A0(reg_out_n3), .A1(reg_out_cipher_sample[121]), 
        .B0(cipher_byte_out[1]), .B1(reg_out_n2), .Y(reg_out_n26) );
  INVX1 reg_out_U300 ( .A(reg_out_n26), .Y(reg_out_n308) );
  AOI22X1 reg_out_U299 ( .A0(reg_out_n4), .A1(reg_out_cipher_sample[120]), 
        .B0(cipher_byte_out[0]), .B1(reg_out_n2), .Y(reg_out_n28) );
  INVX1 reg_out_U298 ( .A(reg_out_n28), .Y(reg_out_n309) );
  AOI22X1 reg_out_U297 ( .A0(reg_out_n3), .A1(reg_out_cipher_sample[127]), 
        .B0(cipher_byte_out[7]), .B1(reg_out_n2), .Y(reg_out_n11) );
  INVX1 reg_out_U296 ( .A(reg_out_n11), .Y(reg_out_n302) );
  AND3X2 reg_out_U295 ( .A(reg_out_rdy1), .B(reg_out_n310), .C(empty), .Y(
        reg_out_n15) );
  AOI22X1 reg_out_U294 ( .A0(reg_out_cipher_sample[103]), .A1(reg_out_n6), 
        .B0(Dout[111]), .B1(reg_out_n282), .Y(reg_out_n38) );
  OAI2BB1X1 reg_out_U293 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[111]), .B0(reg_out_n38), .Y(reg_out_n166) );
  AOI22X1 reg_out_U292 ( .A0(reg_out_cipher_sample[111]), .A1(reg_out_n5), 
        .B0(Dout[119]), .B1(reg_out_n15), .Y(reg_out_n30) );
  OAI2BB1X1 reg_out_U291 ( .A0N(reg_out_cipher_sample[119]), .A1N(reg_out_n298), .B0(reg_out_n30), .Y(reg_out_n158) );
  AOI22X1 reg_out_U290 ( .A0(reg_out_cipher_sample[94]), .A1(reg_out_n7), .B0(
        Dout[102]), .B1(reg_out_n283), .Y(reg_out_n47) );
  OAI2BB1X1 reg_out_U289 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[102]), .B0(reg_out_n47), .Y(reg_out_n175) );
  AOI22X1 reg_out_U288 ( .A0(reg_out_cipher_sample[102]), .A1(reg_out_n6), 
        .B0(Dout[110]), .B1(reg_out_n282), .Y(reg_out_n39) );
  OAI2BB1X1 reg_out_U287 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[110]), .B0(reg_out_n39), .Y(reg_out_n167) );
  AOI22X1 reg_out_U286 ( .A0(reg_out_cipher_sample[93]), .A1(reg_out_n10), 
        .B0(Dout[101]), .B1(reg_out_n283), .Y(reg_out_n48) );
  OAI2BB1X1 reg_out_U285 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[101]), .B0(reg_out_n48), .Y(reg_out_n176) );
  AOI22X1 reg_out_U284 ( .A0(reg_out_cipher_sample[101]), .A1(reg_out_n6), 
        .B0(Dout[109]), .B1(reg_out_n282), .Y(reg_out_n40) );
  OAI2BB1X1 reg_out_U283 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[109]), .B0(reg_out_n40), .Y(reg_out_n168) );
  AOI22X1 reg_out_U282 ( .A0(reg_out_cipher_sample[92]), .A1(reg_out_n7), .B0(
        Dout[100]), .B1(reg_out_n283), .Y(reg_out_n49) );
  OAI2BB1X1 reg_out_U281 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[100]), .B0(reg_out_n49), .Y(reg_out_n177) );
  AOI22X1 reg_out_U280 ( .A0(reg_out_cipher_sample[89]), .A1(reg_out_n7), .B0(
        Dout[97]), .B1(reg_out_n283), .Y(reg_out_n52) );
  OAI2BB1X1 reg_out_U279 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[97]), 
        .B0(reg_out_n52), .Y(reg_out_n180) );
  AOI22X1 reg_out_U278 ( .A0(reg_out_cipher_sample[100]), .A1(reg_out_n6), 
        .B0(Dout[108]), .B1(reg_out_n282), .Y(reg_out_n41) );
  OAI2BB1X1 reg_out_U277 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[108]), .B0(reg_out_n41), .Y(reg_out_n169) );
  AOI22X1 reg_out_U276 ( .A0(reg_out_cipher_sample[98]), .A1(reg_out_n6), .B0(
        Dout[106]), .B1(reg_out_n282), .Y(reg_out_n43) );
  OAI2BB1X1 reg_out_U275 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[106]), .B0(reg_out_n43), .Y(reg_out_n171) );
  AOI22X1 reg_out_U274 ( .A0(reg_out_cipher_sample[97]), .A1(reg_out_n6), .B0(
        Dout[105]), .B1(reg_out_n282), .Y(reg_out_n44) );
  OAI2BB1X1 reg_out_U273 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[105]), .B0(reg_out_n44), .Y(reg_out_n172) );
  AOI22X1 reg_out_U272 ( .A0(reg_out_cipher_sample[96]), .A1(reg_out_n6), .B0(
        Dout[104]), .B1(reg_out_n282), .Y(reg_out_n45) );
  OAI2BB1X1 reg_out_U271 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[104]), .B0(reg_out_n45), .Y(reg_out_n173) );
  AOI22X1 reg_out_U270 ( .A0(reg_out_cipher_sample[39]), .A1(reg_out_n13), 
        .B0(Dout[47]), .B1(reg_out_n287), .Y(reg_out_n102) );
  OAI2BB1X1 reg_out_U269 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[47]), 
        .B0(reg_out_n102), .Y(reg_out_n230) );
  AOI22X1 reg_out_U268 ( .A0(reg_out_cipher_sample[30]), .A1(reg_out_n278), 
        .B0(Dout[38]), .B1(reg_out_n288), .Y(reg_out_n111) );
  OAI2BB1X1 reg_out_U267 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[38]), 
        .B0(reg_out_n111), .Y(reg_out_n239) );
  AOI22X1 reg_out_U266 ( .A0(reg_out_cipher_sample[38]), .A1(reg_out_n13), 
        .B0(Dout[46]), .B1(reg_out_n287), .Y(reg_out_n103) );
  OAI2BB1X1 reg_out_U265 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[46]), 
        .B0(reg_out_n103), .Y(reg_out_n231) );
  AOI22X1 reg_out_U264 ( .A0(reg_out_cipher_sample[29]), .A1(reg_out_n278), 
        .B0(Dout[37]), .B1(reg_out_n288), .Y(reg_out_n112) );
  OAI2BB1X1 reg_out_U263 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[37]), 
        .B0(reg_out_n112), .Y(reg_out_n240) );
  AOI22X1 reg_out_U262 ( .A0(reg_out_cipher_sample[37]), .A1(reg_out_n13), 
        .B0(Dout[45]), .B1(reg_out_n287), .Y(reg_out_n104) );
  OAI2BB1X1 reg_out_U261 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[45]), 
        .B0(reg_out_n104), .Y(reg_out_n232) );
  AOI22X1 reg_out_U260 ( .A0(reg_out_cipher_sample[28]), .A1(reg_out_n278), 
        .B0(Dout[36]), .B1(reg_out_n288), .Y(reg_out_n113) );
  OAI2BB1X1 reg_out_U259 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[36]), 
        .B0(reg_out_n113), .Y(reg_out_n241) );
  AOI22X1 reg_out_U258 ( .A0(reg_out_cipher_sample[36]), .A1(reg_out_n13), 
        .B0(Dout[44]), .B1(reg_out_n287), .Y(reg_out_n105) );
  OAI2BB1X1 reg_out_U257 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[44]), 
        .B0(reg_out_n105), .Y(reg_out_n233) );
  AOI22X1 reg_out_U256 ( .A0(reg_out_cipher_sample[25]), .A1(reg_out_n278), 
        .B0(Dout[33]), .B1(reg_out_n288), .Y(reg_out_n116) );
  OAI2BB1X1 reg_out_U255 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[33]), 
        .B0(reg_out_n116), .Y(reg_out_n244) );
  AOI22X1 reg_out_U254 ( .A0(reg_out_cipher_sample[121]), .A1(reg_out_n4), 
        .B0(Dout[1]), .B1(reg_out_n290), .Y(reg_out_n148) );
  OAI2BB1X1 reg_out_U253 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[1]), 
        .B0(reg_out_n148), .Y(reg_out_n276) );
  AOI22X1 reg_out_U252 ( .A0(reg_out_cipher_sample[0]), .A1(reg_out_n3), .B0(
        Dout[8]), .B1(reg_out_n290), .Y(reg_out_n141) );
  OAI2BB1X1 reg_out_U251 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[8]), 
        .B0(reg_out_n141), .Y(reg_out_n269) );
  AOI22X1 reg_out_U250 ( .A0(reg_out_cipher_sample[119]), .A1(reg_out_n5), 
        .B0(Dout[127]), .B1(reg_out_n15), .Y(reg_out_n14) );
  OAI2BB1X1 reg_out_U249 ( .A0N(reg_out_cipher_sample[127]), .A1N(reg_out_n301), .B0(reg_out_n14), .Y(reg_out_n150) );
  AOI22X1 reg_out_U248 ( .A0(reg_out_cipher_sample[118]), .A1(reg_out_n5), 
        .B0(Dout[126]), .B1(reg_out_n15), .Y(reg_out_n17) );
  OAI2BB1X1 reg_out_U247 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[126]), .B0(reg_out_n17), .Y(reg_out_n151) );
  AOI22X1 reg_out_U246 ( .A0(reg_out_cipher_sample[117]), .A1(reg_out_n5), 
        .B0(Dout[125]), .B1(reg_out_n15), .Y(reg_out_n19) );
  OAI2BB1X1 reg_out_U245 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[125]), .B0(reg_out_n19), .Y(reg_out_n152) );
  AOI22X1 reg_out_U244 ( .A0(reg_out_cipher_sample[95]), .A1(reg_out_n7), .B0(
        Dout[103]), .B1(reg_out_n283), .Y(reg_out_n46) );
  OAI2BB1X1 reg_out_U243 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[103]), .B0(reg_out_n46), .Y(reg_out_n174) );
  AOI22X1 reg_out_U242 ( .A0(reg_out_cipher_sample[62]), .A1(reg_out_n9), .B0(
        Dout[70]), .B1(reg_out_n285), .Y(reg_out_n79) );
  OAI2BB1X1 reg_out_U241 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[70]), 
        .B0(reg_out_n79), .Y(reg_out_n207) );
  AOI22X1 reg_out_U240 ( .A0(reg_out_cipher_sample[70]), .A1(reg_out_n9), .B0(
        Dout[78]), .B1(reg_out_n285), .Y(reg_out_n71) );
  OAI2BB1X1 reg_out_U239 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[78]), 
        .B0(reg_out_n71), .Y(reg_out_n199) );
  AOI22X1 reg_out_U238 ( .A0(reg_out_cipher_sample[110]), .A1(reg_out_n5), 
        .B0(Dout[118]), .B1(reg_out_n15), .Y(reg_out_n31) );
  OAI2BB1X1 reg_out_U237 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[118]), .B0(reg_out_n31), .Y(reg_out_n159) );
  AOI22X1 reg_out_U236 ( .A0(reg_out_cipher_sample[61]), .A1(reg_out_n9), .B0(
        Dout[69]), .B1(reg_out_n285), .Y(reg_out_n80) );
  OAI2BB1X1 reg_out_U235 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[69]), 
        .B0(reg_out_n80), .Y(reg_out_n208) );
  AOI22X1 reg_out_U234 ( .A0(reg_out_cipher_sample[69]), .A1(reg_out_n9), .B0(
        Dout[77]), .B1(reg_out_n285), .Y(reg_out_n72) );
  OAI2BB1X1 reg_out_U233 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[77]), 
        .B0(reg_out_n72), .Y(reg_out_n200) );
  AOI22X1 reg_out_U232 ( .A0(reg_out_cipher_sample[109]), .A1(reg_out_n5), 
        .B0(Dout[117]), .B1(reg_out_n15), .Y(reg_out_n32) );
  OAI2BB1X1 reg_out_U231 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[117]), .B0(reg_out_n32), .Y(reg_out_n160) );
  AOI22X1 reg_out_U230 ( .A0(reg_out_cipher_sample[60]), .A1(reg_out_n9), .B0(
        Dout[68]), .B1(reg_out_n285), .Y(reg_out_n81) );
  OAI2BB1X1 reg_out_U229 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[68]), 
        .B0(reg_out_n81), .Y(reg_out_n209) );
  AOI22X1 reg_out_U228 ( .A0(reg_out_cipher_sample[68]), .A1(reg_out_n9), .B0(
        Dout[76]), .B1(reg_out_n285), .Y(reg_out_n73) );
  OAI2BB1X1 reg_out_U227 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[76]), 
        .B0(reg_out_n73), .Y(reg_out_n201) );
  AOI22X1 reg_out_U226 ( .A0(reg_out_cipher_sample[108]), .A1(reg_out_n5), 
        .B0(Dout[116]), .B1(reg_out_n15), .Y(reg_out_n33) );
  OAI2BB1X1 reg_out_U225 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[116]), .B0(reg_out_n33), .Y(reg_out_n161) );
  AOI22X1 reg_out_U224 ( .A0(reg_out_cipher_sample[59]), .A1(reg_out_n9), .B0(
        Dout[67]), .B1(reg_out_n286), .Y(reg_out_n82) );
  OAI2BB1X1 reg_out_U223 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[67]), 
        .B0(reg_out_n82), .Y(reg_out_n210) );
  AOI22X1 reg_out_U222 ( .A0(reg_out_cipher_sample[67]), .A1(reg_out_n9), .B0(
        Dout[75]), .B1(reg_out_n285), .Y(reg_out_n74) );
  OAI2BB1X1 reg_out_U221 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[75]), 
        .B0(reg_out_n74), .Y(reg_out_n202) );
  AOI22X1 reg_out_U220 ( .A0(reg_out_cipher_sample[91]), .A1(reg_out_n7), .B0(
        Dout[99]), .B1(reg_out_n283), .Y(reg_out_n50) );
  OAI2BB1X1 reg_out_U219 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[99]), 
        .B0(reg_out_n50), .Y(reg_out_n178) );
  AOI22X1 reg_out_U218 ( .A0(reg_out_cipher_sample[58]), .A1(reg_out_n10), 
        .B0(Dout[66]), .B1(reg_out_n286), .Y(reg_out_n83) );
  OAI2BB1X1 reg_out_U217 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[66]), 
        .B0(reg_out_n83), .Y(reg_out_n211) );
  AOI22X1 reg_out_U216 ( .A0(reg_out_cipher_sample[66]), .A1(reg_out_n9), .B0(
        Dout[74]), .B1(reg_out_n285), .Y(reg_out_n75) );
  OAI2BB1X1 reg_out_U215 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[74]), 
        .B0(reg_out_n75), .Y(reg_out_n203) );
  AOI22X1 reg_out_U214 ( .A0(reg_out_cipher_sample[90]), .A1(reg_out_n7), .B0(
        Dout[98]), .B1(reg_out_n283), .Y(reg_out_n51) );
  OAI2BB1X1 reg_out_U213 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[98]), 
        .B0(reg_out_n51), .Y(reg_out_n179) );
  AOI22X1 reg_out_U212 ( .A0(reg_out_cipher_sample[57]), .A1(reg_out_n10), 
        .B0(Dout[65]), .B1(reg_out_n286), .Y(reg_out_n84) );
  OAI2BB1X1 reg_out_U211 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[65]), 
        .B0(reg_out_n84), .Y(reg_out_n212) );
  AOI22X1 reg_out_U210 ( .A0(reg_out_cipher_sample[65]), .A1(reg_out_n9), .B0(
        Dout[73]), .B1(reg_out_n285), .Y(reg_out_n76) );
  OAI2BB1X1 reg_out_U209 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[73]), 
        .B0(reg_out_n76), .Y(reg_out_n204) );
  AOI22X1 reg_out_U208 ( .A0(reg_out_cipher_sample[105]), .A1(reg_out_n6), 
        .B0(Dout[113]), .B1(reg_out_n282), .Y(reg_out_n36) );
  OAI2BB1X1 reg_out_U207 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[113]), .B0(reg_out_n36), .Y(reg_out_n164) );
  AOI22X1 reg_out_U206 ( .A0(reg_out_cipher_sample[56]), .A1(reg_out_n10), 
        .B0(Dout[64]), .B1(reg_out_n286), .Y(reg_out_n85) );
  OAI2BB1X1 reg_out_U205 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[64]), 
        .B0(reg_out_n85), .Y(reg_out_n213) );
  AOI22X1 reg_out_U204 ( .A0(reg_out_cipher_sample[64]), .A1(reg_out_n9), .B0(
        Dout[72]), .B1(reg_out_n285), .Y(reg_out_n77) );
  OAI2BB1X1 reg_out_U203 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[72]), 
        .B0(reg_out_n77), .Y(reg_out_n205) );
  AOI22X1 reg_out_U202 ( .A0(reg_out_cipher_sample[99]), .A1(reg_out_n6), .B0(
        Dout[107]), .B1(reg_out_n282), .Y(reg_out_n42) );
  OAI2BB1X1 reg_out_U201 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[107]), .B0(reg_out_n42), .Y(reg_out_n170) );
  AOI22X1 reg_out_U200 ( .A0(reg_out_cipher_sample[27]), .A1(reg_out_n278), 
        .B0(Dout[35]), .B1(reg_out_n288), .Y(reg_out_n114) );
  OAI2BB1X1 reg_out_U199 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[35]), 
        .B0(reg_out_n114), .Y(reg_out_n242) );
  AOI22X1 reg_out_U198 ( .A0(reg_out_cipher_sample[26]), .A1(reg_out_n278), 
        .B0(Dout[34]), .B1(reg_out_n288), .Y(reg_out_n115) );
  OAI2BB1X1 reg_out_U197 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[34]), 
        .B0(reg_out_n115), .Y(reg_out_n243) );
  AOI22X1 reg_out_U196 ( .A0(reg_out_cipher_sample[24]), .A1(reg_out_n278), 
        .B0(Dout[32]), .B1(reg_out_n288), .Y(reg_out_n117) );
  OAI2BB1X1 reg_out_U195 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[32]), 
        .B0(reg_out_n117), .Y(reg_out_n245) );
  AOI22X1 reg_out_U194 ( .A0(reg_out_cipher_sample[123]), .A1(reg_out_n4), 
        .B0(Dout[3]), .B1(reg_out_n290), .Y(reg_out_n146) );
  OAI2BB1X1 reg_out_U193 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[3]), 
        .B0(reg_out_n146), .Y(reg_out_n274) );
  AOI22X1 reg_out_U192 ( .A0(reg_out_cipher_sample[122]), .A1(reg_out_n4), 
        .B0(Dout[2]), .B1(reg_out_n290), .Y(reg_out_n147) );
  OAI2BB1X1 reg_out_U191 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[2]), 
        .B0(reg_out_n147), .Y(reg_out_n275) );
  AOI22X1 reg_out_U190 ( .A0(reg_out_cipher_sample[2]), .A1(reg_out_n3), .B0(
        Dout[10]), .B1(reg_out_n290), .Y(reg_out_n139) );
  OAI2BB1X1 reg_out_U189 ( .A0N(reg_out_n292), .A1N(reg_out_cipher_sample[10]), 
        .B0(reg_out_n139), .Y(reg_out_n267) );
  AOI22X1 reg_out_U188 ( .A0(reg_out_cipher_sample[120]), .A1(reg_out_n4), 
        .B0(Dout[0]), .B1(reg_out_n290), .Y(reg_out_n149) );
  OAI2BB1X1 reg_out_U187 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[0]), 
        .B0(reg_out_n149), .Y(reg_out_n277) );
  AOI22X1 reg_out_U186 ( .A0(reg_out_cipher_sample[116]), .A1(reg_out_n5), 
        .B0(Dout[124]), .B1(reg_out_n15), .Y(reg_out_n21) );
  OAI2BB1X1 reg_out_U185 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[124]), .B0(reg_out_n21), .Y(reg_out_n153) );
  AOI22X1 reg_out_U184 ( .A0(reg_out_cipher_sample[114]), .A1(reg_out_n5), 
        .B0(Dout[122]), .B1(reg_out_n15), .Y(reg_out_n25) );
  OAI2BB1X1 reg_out_U183 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[122]), .B0(reg_out_n25), .Y(reg_out_n155) );
  AOI22X1 reg_out_U182 ( .A0(reg_out_cipher_sample[113]), .A1(reg_out_n5), 
        .B0(Dout[121]), .B1(reg_out_n15), .Y(reg_out_n27) );
  OAI2BB1X1 reg_out_U181 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[121]), .B0(reg_out_n27), .Y(reg_out_n156) );
  AOI22X1 reg_out_U180 ( .A0(reg_out_cipher_sample[112]), .A1(reg_out_n5), 
        .B0(Dout[120]), .B1(reg_out_n15), .Y(reg_out_n29) );
  OAI2BB1X1 reg_out_U179 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[120]), .B0(reg_out_n29), .Y(reg_out_n157) );
  AOI22X1 reg_out_U178 ( .A0(reg_out_cipher_sample[107]), .A1(reg_out_n6), 
        .B0(Dout[115]), .B1(reg_out_n282), .Y(reg_out_n34) );
  OAI2BB1X1 reg_out_U177 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[115]), .B0(reg_out_n34), .Y(reg_out_n162) );
  AOI22X1 reg_out_U176 ( .A0(reg_out_cipher_sample[106]), .A1(reg_out_n6), 
        .B0(Dout[114]), .B1(reg_out_n282), .Y(reg_out_n35) );
  OAI2BB1X1 reg_out_U175 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[114]), .B0(reg_out_n35), .Y(reg_out_n163) );
  AOI22X1 reg_out_U174 ( .A0(reg_out_cipher_sample[88]), .A1(reg_out_n7), .B0(
        Dout[96]), .B1(reg_out_n283), .Y(reg_out_n53) );
  OAI2BB1X1 reg_out_U173 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[96]), 
        .B0(reg_out_n53), .Y(reg_out_n181) );
  AOI22X1 reg_out_U172 ( .A0(reg_out_cipher_sample[104]), .A1(reg_out_n6), 
        .B0(Dout[112]), .B1(reg_out_n282), .Y(reg_out_n37) );
  OAI2BB1X1 reg_out_U171 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[112]), .B0(reg_out_n37), .Y(reg_out_n165) );
  AOI22X1 reg_out_U170 ( .A0(reg_out_cipher_sample[47]), .A1(reg_out_n13), 
        .B0(Dout[55]), .B1(reg_out_n287), .Y(reg_out_n94) );
  OAI2BB1X1 reg_out_U169 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[55]), 
        .B0(reg_out_n94), .Y(reg_out_n222) );
  AOI22X1 reg_out_U168 ( .A0(reg_out_cipher_sample[46]), .A1(reg_out_n13), 
        .B0(Dout[54]), .B1(reg_out_n287), .Y(reg_out_n95) );
  OAI2BB1X1 reg_out_U167 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[54]), 
        .B0(reg_out_n95), .Y(reg_out_n223) );
  AOI22X1 reg_out_U166 ( .A0(reg_out_cipher_sample[45]), .A1(reg_out_n13), 
        .B0(Dout[53]), .B1(reg_out_n287), .Y(reg_out_n96) );
  OAI2BB1X1 reg_out_U165 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[53]), 
        .B0(reg_out_n96), .Y(reg_out_n224) );
  AOI22X1 reg_out_U164 ( .A0(reg_out_cipher_sample[44]), .A1(reg_out_n13), 
        .B0(Dout[52]), .B1(reg_out_n287), .Y(reg_out_n97) );
  OAI2BB1X1 reg_out_U163 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[52]), 
        .B0(reg_out_n97), .Y(reg_out_n225) );
  AOI22X1 reg_out_U162 ( .A0(reg_out_cipher_sample[33]), .A1(reg_out_n278), 
        .B0(Dout[41]), .B1(reg_out_n288), .Y(reg_out_n108) );
  OAI2BB1X1 reg_out_U161 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[41]), 
        .B0(reg_out_n108), .Y(reg_out_n236) );
  AOI22X1 reg_out_U160 ( .A0(reg_out_cipher_sample[41]), .A1(reg_out_n13), 
        .B0(Dout[49]), .B1(reg_out_n287), .Y(reg_out_n100) );
  OAI2BB1X1 reg_out_U159 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[49]), 
        .B0(reg_out_n100), .Y(reg_out_n228) );
  AOI22X1 reg_out_U158 ( .A0(reg_out_cipher_sample[7]), .A1(reg_out_n3), .B0(
        Dout[15]), .B1(reg_out_n15), .Y(reg_out_n134) );
  OAI2BB1X1 reg_out_U157 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[15]), 
        .B0(reg_out_n134), .Y(reg_out_n262) );
  AOI22X1 reg_out_U156 ( .A0(reg_out_cipher_sample[15]), .A1(reg_out_n279), 
        .B0(Dout[23]), .B1(reg_out_n289), .Y(reg_out_n126) );
  OAI2BB1X1 reg_out_U155 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[23]), 
        .B0(reg_out_n126), .Y(reg_out_n254) );
  AOI22X1 reg_out_U154 ( .A0(reg_out_cipher_sample[126]), .A1(reg_out_n4), 
        .B0(Dout[6]), .B1(reg_out_n290), .Y(reg_out_n143) );
  OAI2BB1X1 reg_out_U153 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[6]), 
        .B0(reg_out_n143), .Y(reg_out_n271) );
  AOI22X1 reg_out_U152 ( .A0(reg_out_cipher_sample[6]), .A1(reg_out_n3), .B0(
        Dout[14]), .B1(reg_out_n15), .Y(reg_out_n135) );
  OAI2BB1X1 reg_out_U151 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[14]), 
        .B0(reg_out_n135), .Y(reg_out_n263) );
  AOI22X1 reg_out_U150 ( .A0(reg_out_cipher_sample[14]), .A1(reg_out_n279), 
        .B0(Dout[22]), .B1(reg_out_n289), .Y(reg_out_n127) );
  OAI2BB1X1 reg_out_U149 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[22]), 
        .B0(reg_out_n127), .Y(reg_out_n255) );
  AOI22X1 reg_out_U148 ( .A0(reg_out_cipher_sample[125]), .A1(reg_out_n4), 
        .B0(Dout[5]), .B1(reg_out_n290), .Y(reg_out_n144) );
  OAI2BB1X1 reg_out_U147 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[5]), 
        .B0(reg_out_n144), .Y(reg_out_n272) );
  AOI22X1 reg_out_U146 ( .A0(reg_out_cipher_sample[5]), .A1(reg_out_n3), .B0(
        Dout[13]), .B1(reg_out_n15), .Y(reg_out_n136) );
  OAI2BB1X1 reg_out_U145 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[13]), 
        .B0(reg_out_n136), .Y(reg_out_n264) );
  AOI22X1 reg_out_U144 ( .A0(reg_out_cipher_sample[13]), .A1(reg_out_n279), 
        .B0(Dout[21]), .B1(reg_out_n289), .Y(reg_out_n128) );
  OAI2BB1X1 reg_out_U143 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[21]), 
        .B0(reg_out_n128), .Y(reg_out_n256) );
  AOI22X1 reg_out_U142 ( .A0(reg_out_cipher_sample[124]), .A1(reg_out_n4), 
        .B0(Dout[4]), .B1(reg_out_n290), .Y(reg_out_n145) );
  OAI2BB1X1 reg_out_U141 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[4]), 
        .B0(reg_out_n145), .Y(reg_out_n273) );
  AOI22X1 reg_out_U140 ( .A0(reg_out_cipher_sample[12]), .A1(reg_out_n279), 
        .B0(Dout[20]), .B1(reg_out_n289), .Y(reg_out_n129) );
  OAI2BB1X1 reg_out_U139 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[20]), 
        .B0(reg_out_n129), .Y(reg_out_n257) );
  AOI22X1 reg_out_U138 ( .A0(reg_out_cipher_sample[1]), .A1(reg_out_n3), .B0(
        Dout[9]), .B1(reg_out_n15), .Y(reg_out_n140) );
  OAI2BB1X1 reg_out_U137 ( .A0N(reg_out_n294), .A1N(reg_out_cipher_sample[9]), 
        .B0(reg_out_n140), .Y(reg_out_n268) );
  AOI22X1 reg_out_U136 ( .A0(reg_out_cipher_sample[9]), .A1(reg_out_n3), .B0(
        Dout[17]), .B1(reg_out_n15), .Y(reg_out_n132) );
  OAI2BB1X1 reg_out_U135 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[17]), 
        .B0(reg_out_n132), .Y(reg_out_n260) );
  AOI22X1 reg_out_U134 ( .A0(reg_out_cipher_sample[86]), .A1(reg_out_n7), .B0(
        Dout[94]), .B1(reg_out_n283), .Y(reg_out_n55) );
  OAI2BB1X1 reg_out_U133 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[94]), 
        .B0(reg_out_n55), .Y(reg_out_n183) );
  AOI22X1 reg_out_U132 ( .A0(reg_out_cipher_sample[85]), .A1(reg_out_n7), .B0(
        Dout[93]), .B1(reg_out_n283), .Y(reg_out_n56) );
  OAI2BB1X1 reg_out_U131 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[93]), 
        .B0(reg_out_n56), .Y(reg_out_n184) );
  AOI22X1 reg_out_U130 ( .A0(reg_out_cipher_sample[84]), .A1(reg_out_n7), .B0(
        Dout[92]), .B1(reg_out_n283), .Y(reg_out_n57) );
  OAI2BB1X1 reg_out_U129 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[92]), 
        .B0(reg_out_n57), .Y(reg_out_n185) );
  AOI22X1 reg_out_U128 ( .A0(reg_out_cipher_sample[71]), .A1(reg_out_n8), .B0(
        Dout[79]), .B1(reg_out_n285), .Y(reg_out_n70) );
  OAI2BB1X1 reg_out_U127 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[79]), 
        .B0(reg_out_n70), .Y(reg_out_n198) );
  AOI22X1 reg_out_U126 ( .A0(reg_out_cipher_sample[79]), .A1(reg_out_n8), .B0(
        Dout[87]), .B1(reg_out_n284), .Y(reg_out_n62) );
  OAI2BB1X1 reg_out_U125 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[87]), 
        .B0(reg_out_n62), .Y(reg_out_n190) );
  AOI22X1 reg_out_U124 ( .A0(reg_out_cipher_sample[78]), .A1(reg_out_n8), .B0(
        Dout[86]), .B1(reg_out_n284), .Y(reg_out_n63) );
  OAI2BB1X1 reg_out_U123 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[86]), 
        .B0(reg_out_n63), .Y(reg_out_n191) );
  AOI22X1 reg_out_U122 ( .A0(reg_out_cipher_sample[77]), .A1(reg_out_n8), .B0(
        Dout[85]), .B1(reg_out_n284), .Y(reg_out_n64) );
  OAI2BB1X1 reg_out_U121 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[85]), 
        .B0(reg_out_n64), .Y(reg_out_n192) );
  AOI22X1 reg_out_U120 ( .A0(reg_out_cipher_sample[76]), .A1(reg_out_n8), .B0(
        Dout[84]), .B1(reg_out_n284), .Y(reg_out_n65) );
  OAI2BB1X1 reg_out_U119 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[84]), 
        .B0(reg_out_n65), .Y(reg_out_n193) );
  AOI22X1 reg_out_U118 ( .A0(reg_out_cipher_sample[75]), .A1(reg_out_n8), .B0(
        Dout[83]), .B1(reg_out_n284), .Y(reg_out_n66) );
  OAI2BB1X1 reg_out_U117 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[83]), 
        .B0(reg_out_n66), .Y(reg_out_n194) );
  AOI22X1 reg_out_U116 ( .A0(reg_out_cipher_sample[74]), .A1(reg_out_n8), .B0(
        Dout[82]), .B1(reg_out_n284), .Y(reg_out_n67) );
  OAI2BB1X1 reg_out_U115 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[82]), 
        .B0(reg_out_n67), .Y(reg_out_n195) );
  AOI22X1 reg_out_U114 ( .A0(reg_out_cipher_sample[73]), .A1(reg_out_n8), .B0(
        Dout[81]), .B1(reg_out_n284), .Y(reg_out_n68) );
  OAI2BB1X1 reg_out_U113 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[81]), 
        .B0(reg_out_n68), .Y(reg_out_n196) );
  AOI22X1 reg_out_U112 ( .A0(reg_out_cipher_sample[72]), .A1(reg_out_n8), .B0(
        Dout[80]), .B1(reg_out_n284), .Y(reg_out_n69) );
  OAI2BB1X1 reg_out_U111 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[80]), 
        .B0(reg_out_n69), .Y(reg_out_n197) );
  AOI22X1 reg_out_U110 ( .A0(reg_out_cipher_sample[3]), .A1(reg_out_n3), .B0(
        Dout[11]), .B1(reg_out_n15), .Y(reg_out_n138) );
  OAI2BB1X1 reg_out_U109 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[11]), 
        .B0(reg_out_n138), .Y(reg_out_n266) );
  AOI22X1 reg_out_U108 ( .A0(reg_out_cipher_sample[115]), .A1(reg_out_n5), 
        .B0(Dout[123]), .B1(reg_out_n15), .Y(reg_out_n23) );
  OAI2BB1X1 reg_out_U107 ( .A0N(reg_out_n293), .A1N(reg_out_cipher_sample[123]), .B0(reg_out_n23), .Y(reg_out_n154) );
  AOI22X1 reg_out_U106 ( .A0(reg_out_cipher_sample[35]), .A1(reg_out_n278), 
        .B0(Dout[43]), .B1(reg_out_n288), .Y(reg_out_n106) );
  OAI2BB1X1 reg_out_U105 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[43]), 
        .B0(reg_out_n106), .Y(reg_out_n234) );
  AOI22X1 reg_out_U104 ( .A0(reg_out_cipher_sample[43]), .A1(reg_out_n13), 
        .B0(Dout[51]), .B1(reg_out_n287), .Y(reg_out_n98) );
  OAI2BB1X1 reg_out_U103 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[51]), 
        .B0(reg_out_n98), .Y(reg_out_n226) );
  AOI22X1 reg_out_U102 ( .A0(reg_out_cipher_sample[34]), .A1(reg_out_n278), 
        .B0(Dout[42]), .B1(reg_out_n288), .Y(reg_out_n107) );
  OAI2BB1X1 reg_out_U101 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[42]), 
        .B0(reg_out_n107), .Y(reg_out_n235) );
  AOI22X1 reg_out_U100 ( .A0(reg_out_cipher_sample[42]), .A1(reg_out_n13), 
        .B0(Dout[50]), .B1(reg_out_n287), .Y(reg_out_n99) );
  OAI2BB1X1 reg_out_U99 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[50]), 
        .B0(reg_out_n99), .Y(reg_out_n227) );
  AOI22X1 reg_out_U98 ( .A0(reg_out_cipher_sample[32]), .A1(reg_out_n278), 
        .B0(Dout[40]), .B1(reg_out_n288), .Y(reg_out_n109) );
  OAI2BB1X1 reg_out_U97 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[40]), 
        .B0(reg_out_n109), .Y(reg_out_n237) );
  AOI22X1 reg_out_U96 ( .A0(reg_out_cipher_sample[40]), .A1(reg_out_n13), .B0(
        Dout[48]), .B1(reg_out_n287), .Y(reg_out_n101) );
  OAI2BB1X1 reg_out_U95 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[48]), 
        .B0(reg_out_n101), .Y(reg_out_n229) );
  AOI22X1 reg_out_U94 ( .A0(reg_out_cipher_sample[4]), .A1(reg_out_n280), .B0(
        Dout[12]), .B1(reg_out_n15), .Y(reg_out_n137) );
  OAI2BB1X1 reg_out_U93 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[12]), 
        .B0(reg_out_n137), .Y(reg_out_n265) );
  AOI22X1 reg_out_U92 ( .A0(reg_out_cipher_sample[11]), .A1(reg_out_n4), .B0(
        Dout[19]), .B1(reg_out_n15), .Y(reg_out_n130) );
  OAI2BB1X1 reg_out_U91 ( .A0N(reg_out_n299), .A1N(reg_out_cipher_sample[19]), 
        .B0(reg_out_n130), .Y(reg_out_n258) );
  AOI22X1 reg_out_U90 ( .A0(reg_out_cipher_sample[10]), .A1(reg_out_n4), .B0(
        Dout[18]), .B1(reg_out_n15), .Y(reg_out_n131) );
  OAI2BB1X1 reg_out_U89 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[18]), 
        .B0(reg_out_n131), .Y(reg_out_n259) );
  AOI22X1 reg_out_U88 ( .A0(reg_out_cipher_sample[8]), .A1(reg_out_n280), .B0(
        Dout[16]), .B1(reg_out_n15), .Y(reg_out_n133) );
  OAI2BB1X1 reg_out_U87 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[16]), 
        .B0(reg_out_n133), .Y(reg_out_n261) );
  AOI22X1 reg_out_U86 ( .A0(reg_out_cipher_sample[83]), .A1(reg_out_n7), .B0(
        Dout[91]), .B1(reg_out_n284), .Y(reg_out_n58) );
  OAI2BB1X1 reg_out_U85 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[91]), 
        .B0(reg_out_n58), .Y(reg_out_n186) );
  AOI22X1 reg_out_U84 ( .A0(reg_out_cipher_sample[82]), .A1(reg_out_n8), .B0(
        Dout[90]), .B1(reg_out_n284), .Y(reg_out_n59) );
  OAI2BB1X1 reg_out_U83 ( .A0N(reg_out_n295), .A1N(reg_out_cipher_sample[90]), 
        .B0(reg_out_n59), .Y(reg_out_n187) );
  AOI22X1 reg_out_U82 ( .A0(reg_out_cipher_sample[81]), .A1(reg_out_n8), .B0(
        Dout[89]), .B1(reg_out_n284), .Y(reg_out_n60) );
  OAI2BB1X1 reg_out_U81 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[89]), 
        .B0(reg_out_n60), .Y(reg_out_n188) );
  AOI22X1 reg_out_U80 ( .A0(reg_out_cipher_sample[80]), .A1(reg_out_n8), .B0(
        Dout[88]), .B1(reg_out_n284), .Y(reg_out_n61) );
  OAI2BB1X1 reg_out_U79 ( .A0N(reg_out_n296), .A1N(reg_out_cipher_sample[88]), 
        .B0(reg_out_n61), .Y(reg_out_n189) );
  AOI22X1 reg_out_U78 ( .A0(reg_out_cipher_sample[55]), .A1(reg_out_n10), .B0(
        Dout[63]), .B1(reg_out_n286), .Y(reg_out_n86) );
  OAI2BB1X1 reg_out_U77 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[63]), 
        .B0(reg_out_n86), .Y(reg_out_n214) );
  AOI22X1 reg_out_U76 ( .A0(reg_out_cipher_sample[54]), .A1(reg_out_n10), .B0(
        Dout[62]), .B1(reg_out_n286), .Y(reg_out_n87) );
  OAI2BB1X1 reg_out_U75 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[62]), 
        .B0(reg_out_n87), .Y(reg_out_n215) );
  AOI22X1 reg_out_U74 ( .A0(reg_out_cipher_sample[53]), .A1(reg_out_n10), .B0(
        Dout[61]), .B1(reg_out_n286), .Y(reg_out_n88) );
  OAI2BB1X1 reg_out_U73 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[61]), 
        .B0(reg_out_n88), .Y(reg_out_n216) );
  AOI22X1 reg_out_U72 ( .A0(reg_out_cipher_sample[52]), .A1(reg_out_n10), .B0(
        Dout[60]), .B1(reg_out_n286), .Y(reg_out_n89) );
  OAI2BB1X1 reg_out_U71 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[60]), 
        .B0(reg_out_n89), .Y(reg_out_n217) );
  AOI22X1 reg_out_U70 ( .A0(reg_out_cipher_sample[49]), .A1(reg_out_n10), .B0(
        Dout[57]), .B1(reg_out_n286), .Y(reg_out_n92) );
  OAI2BB1X1 reg_out_U69 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[57]), 
        .B0(reg_out_n92), .Y(reg_out_n220) );
  AOI22X1 reg_out_U68 ( .A0(reg_out_cipher_sample[23]), .A1(reg_out_n279), 
        .B0(Dout[31]), .B1(reg_out_n289), .Y(reg_out_n118) );
  OAI2BB1X1 reg_out_U67 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[31]), 
        .B0(reg_out_n118), .Y(reg_out_n246) );
  AOI22X1 reg_out_U66 ( .A0(reg_out_cipher_sample[22]), .A1(reg_out_n279), 
        .B0(Dout[30]), .B1(reg_out_n289), .Y(reg_out_n119) );
  OAI2BB1X1 reg_out_U65 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[30]), 
        .B0(reg_out_n119), .Y(reg_out_n247) );
  AOI22X1 reg_out_U64 ( .A0(reg_out_cipher_sample[21]), .A1(reg_out_n279), 
        .B0(Dout[29]), .B1(reg_out_n289), .Y(reg_out_n120) );
  OAI2BB1X1 reg_out_U63 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[29]), 
        .B0(reg_out_n120), .Y(reg_out_n248) );
  AOI22X1 reg_out_U62 ( .A0(reg_out_cipher_sample[31]), .A1(reg_out_n278), 
        .B0(Dout[39]), .B1(reg_out_n288), .Y(reg_out_n110) );
  OAI2BB1X1 reg_out_U61 ( .A0N(reg_out_n300), .A1N(reg_out_cipher_sample[39]), 
        .B0(reg_out_n110), .Y(reg_out_n238) );
  AOI22X1 reg_out_U60 ( .A0(reg_out_cipher_sample[87]), .A1(reg_out_n7), .B0(
        Dout[95]), .B1(reg_out_n283), .Y(reg_out_n54) );
  OAI2BB1X1 reg_out_U59 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[95]), 
        .B0(reg_out_n54), .Y(reg_out_n182) );
  AOI22X1 reg_out_U58 ( .A0(reg_out_cipher_sample[63]), .A1(reg_out_n9), .B0(
        Dout[71]), .B1(reg_out_n285), .Y(reg_out_n78) );
  OAI2BB1X1 reg_out_U57 ( .A0N(reg_out_n297), .A1N(reg_out_cipher_sample[71]), 
        .B0(reg_out_n78), .Y(reg_out_n206) );
  AOI22X1 reg_out_U56 ( .A0(reg_out_cipher_sample[51]), .A1(reg_out_n10), .B0(
        Dout[59]), .B1(reg_out_n286), .Y(reg_out_n90) );
  OAI2BB1X1 reg_out_U55 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[59]), 
        .B0(reg_out_n90), .Y(reg_out_n218) );
  AOI22X1 reg_out_U54 ( .A0(reg_out_cipher_sample[50]), .A1(reg_out_n10), .B0(
        Dout[58]), .B1(reg_out_n286), .Y(reg_out_n91) );
  OAI2BB1X1 reg_out_U53 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[58]), 
        .B0(reg_out_n91), .Y(reg_out_n219) );
  AOI22X1 reg_out_U52 ( .A0(reg_out_cipher_sample[48]), .A1(reg_out_n10), .B0(
        Dout[56]), .B1(reg_out_n286), .Y(reg_out_n93) );
  OAI2BB1X1 reg_out_U51 ( .A0N(reg_out_n298), .A1N(reg_out_cipher_sample[56]), 
        .B0(reg_out_n93), .Y(reg_out_n221) );
  AOI22X1 reg_out_U50 ( .A0(reg_out_cipher_sample[20]), .A1(reg_out_n279), 
        .B0(Dout[28]), .B1(reg_out_n289), .Y(reg_out_n121) );
  OAI2BB1X1 reg_out_U49 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[28]), 
        .B0(reg_out_n121), .Y(reg_out_n249) );
  AOI22X1 reg_out_U48 ( .A0(reg_out_cipher_sample[18]), .A1(reg_out_n279), 
        .B0(Dout[26]), .B1(reg_out_n289), .Y(reg_out_n123) );
  OAI2BB1X1 reg_out_U47 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[26]), 
        .B0(reg_out_n123), .Y(reg_out_n251) );
  AOI22X1 reg_out_U46 ( .A0(reg_out_cipher_sample[17]), .A1(reg_out_n279), 
        .B0(Dout[25]), .B1(reg_out_n289), .Y(reg_out_n124) );
  OAI2BB1X1 reg_out_U45 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[25]), 
        .B0(reg_out_n124), .Y(reg_out_n252) );
  AOI22X1 reg_out_U44 ( .A0(reg_out_cipher_sample[16]), .A1(reg_out_n279), 
        .B0(Dout[24]), .B1(reg_out_n289), .Y(reg_out_n125) );
  OAI2BB1X1 reg_out_U43 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[24]), 
        .B0(reg_out_n125), .Y(reg_out_n253) );
  AOI22X1 reg_out_U42 ( .A0(reg_out_cipher_sample[127]), .A1(reg_out_n4), .B0(
        Dout[7]), .B1(reg_out_n290), .Y(reg_out_n142) );
  OAI2BB1X1 reg_out_U41 ( .A0N(reg_out_n292), .A1N(reg_out_cipher_sample[7]), 
        .B0(reg_out_n142), .Y(reg_out_n270) );
  AOI22X1 reg_out_U40 ( .A0(reg_out_cipher_sample[19]), .A1(reg_out_n279), 
        .B0(Dout[27]), .B1(reg_out_n289), .Y(reg_out_n122) );
  OAI2BB1X1 reg_out_U39 ( .A0N(reg_out_n301), .A1N(reg_out_cipher_sample[27]), 
        .B0(reg_out_n122), .Y(reg_out_n250) );
  NAND3BX1 reg_out_U38 ( .AN(empty), .B(reg_out_n310), .C(reg_out_rdy1), .Y(
        reg_out_n12) );
  BUFX3 reg_out_U37 ( .A(reg_out_n12), .Y(reg_out_n2) );
  INVX1 reg_out_U36 ( .A(reg_out_n15), .Y(reg_out_n291) );
  INVX1 reg_out_U35 ( .A(reg_out_n291), .Y(reg_out_n289) );
  INVX1 reg_out_U34 ( .A(reg_out_n291), .Y(reg_out_n288) );
  INVX1 reg_out_U33 ( .A(reg_out_n291), .Y(reg_out_n287) );
  INVX1 reg_out_U32 ( .A(reg_out_n291), .Y(reg_out_n286) );
  INVX1 reg_out_U31 ( .A(reg_out_n291), .Y(reg_out_n285) );
  INVX1 reg_out_U30 ( .A(reg_out_n291), .Y(reg_out_n284) );
  INVX1 reg_out_U29 ( .A(reg_out_n291), .Y(reg_out_n283) );
  INVX1 reg_out_U28 ( .A(reg_out_n291), .Y(reg_out_n282) );
  INVX1 reg_out_U27 ( .A(reg_out_n2), .Y(reg_out_n4) );
  INVX1 reg_out_U26 ( .A(reg_out_n291), .Y(reg_out_n290) );
  INVX1 reg_out_U25 ( .A(reg_out_n2), .Y(reg_out_n3) );
  INVX1 reg_out_U24 ( .A(reg_out_n4), .Y(reg_out_n281) );
  OR2X2 reg_out_U23 ( .A(reg_out_n290), .B(reg_out_n280), .Y(reg_out_n1) );
  INVX1 reg_out_U22 ( .A(reg_out_n2), .Y(reg_out_n279) );
  INVX1 reg_out_U21 ( .A(reg_out_n2), .Y(reg_out_n278) );
  INVX1 reg_out_U20 ( .A(reg_out_n2), .Y(reg_out_n13) );
  INVX1 reg_out_U19 ( .A(reg_out_n281), .Y(reg_out_n10) );
  INVX1 reg_out_U18 ( .A(reg_out_n281), .Y(reg_out_n9) );
  INVX1 reg_out_U17 ( .A(reg_out_n281), .Y(reg_out_n8) );
  INVX1 reg_out_U16 ( .A(reg_out_n281), .Y(reg_out_n7) );
  INVX1 reg_out_U15 ( .A(reg_out_n281), .Y(reg_out_n6) );
  INVX1 reg_out_U14 ( .A(reg_out_n281), .Y(reg_out_n5) );
  INVX1 reg_out_U13 ( .A(reg_out_n1), .Y(reg_out_n292) );
  INVX1 reg_out_U12 ( .A(reg_out_n2), .Y(reg_out_n280) );
  INVX1 reg_out_U11 ( .A(reg_out_n1), .Y(reg_out_n293) );
  INVX1 reg_out_U10 ( .A(reg_out_n1), .Y(reg_out_n301) );
  INVX1 reg_out_U9 ( .A(reg_out_n1), .Y(reg_out_n300) );
  INVX1 reg_out_U8 ( .A(reg_out_n1), .Y(reg_out_n299) );
  INVX1 reg_out_U7 ( .A(reg_out_n1), .Y(reg_out_n298) );
  INVX1 reg_out_U6 ( .A(reg_out_n1), .Y(reg_out_n297) );
  INVX1 reg_out_U5 ( .A(reg_out_n1), .Y(reg_out_n296) );
  INVX1 reg_out_U4 ( .A(reg_out_n1), .Y(reg_out_n294) );
  INVX1 reg_out_U3 ( .A(reg_out_n1), .Y(reg_out_n295) );
  DFFRHQX1 reg_out_rdy2_reg ( .D(reg_out_rdy1), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(reg_out_rdy2) );
  DFFRHQX1 reg_out_rdy0_reg ( .D(ready), .CK(clk_48Mhz), .RN(reset_n), .Q(
        reg_out_rdy0) );
  DFFRHQX1 reg_out_rdy1_reg ( .D(reg_out_rdy0), .CK(clk_48Mhz), .RN(reset_n), 
        .Q(reg_out_rdy1) );
  DFFRHQX1 reg_out_cipher_byte_reg_0_ ( .D(reg_out_n309), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[0]) );
  DFFRHQX1 reg_out_cipher_byte_reg_1_ ( .D(reg_out_n308), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[1]) );
  DFFRHQX1 reg_out_cipher_byte_reg_2_ ( .D(reg_out_n307), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[2]) );
  DFFRHQX1 reg_out_cipher_byte_reg_3_ ( .D(reg_out_n306), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[3]) );
  DFFRHQX1 reg_out_cipher_byte_reg_4_ ( .D(reg_out_n305), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[4]) );
  DFFRHQX1 reg_out_cipher_byte_reg_5_ ( .D(reg_out_n304), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[5]) );
  DFFRHQX1 reg_out_cipher_byte_reg_6_ ( .D(reg_out_n303), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[6]) );
  DFFRHQX1 reg_out_cipher_byte_reg_7_ ( .D(reg_out_n302), .CK(clk_48Mhz), .RN(
        reset_n), .Q(cipher_byte_out[7]) );
  DFFRHQX1 reg_out_cipher_sample_reg_127_ ( .D(reg_out_n150), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[127]) );
  DFFRHQX1 reg_out_cipher_sample_reg_120_ ( .D(reg_out_n157), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[120]) );
  DFFRHQX1 reg_out_cipher_sample_reg_121_ ( .D(reg_out_n156), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[121]) );
  DFFRHQX1 reg_out_cipher_sample_reg_122_ ( .D(reg_out_n155), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[122]) );
  DFFRHQX1 reg_out_cipher_sample_reg_123_ ( .D(reg_out_n154), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[123]) );
  DFFRHQX1 reg_out_cipher_sample_reg_124_ ( .D(reg_out_n153), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[124]) );
  DFFRHQX1 reg_out_cipher_sample_reg_125_ ( .D(reg_out_n152), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[125]) );
  DFFRHQX1 reg_out_cipher_sample_reg_126_ ( .D(reg_out_n151), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[126]) );
  DFFRHQX1 reg_out_cipher_sample_reg_119_ ( .D(reg_out_n158), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[119]) );
  DFFRHQX1 reg_out_cipher_sample_reg_112_ ( .D(reg_out_n165), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[112]) );
  DFFRHQX1 reg_out_cipher_sample_reg_104_ ( .D(reg_out_n173), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[104]) );
  DFFRHQX1 reg_out_cipher_sample_reg_96_ ( .D(reg_out_n181), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[96]) );
  DFFRHQX1 reg_out_cipher_sample_reg_88_ ( .D(reg_out_n189), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[88]) );
  DFFRHQX1 reg_out_cipher_sample_reg_80_ ( .D(reg_out_n197), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[80]) );
  DFFRHQX1 reg_out_cipher_sample_reg_72_ ( .D(reg_out_n205), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[72]) );
  DFFRHQX1 reg_out_cipher_sample_reg_64_ ( .D(reg_out_n213), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[64]) );
  DFFRHQX1 reg_out_cipher_sample_reg_56_ ( .D(reg_out_n221), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[56]) );
  DFFRHQX1 reg_out_cipher_sample_reg_48_ ( .D(reg_out_n229), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[48]) );
  DFFRHQX1 reg_out_cipher_sample_reg_40_ ( .D(reg_out_n237), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[40]) );
  DFFRHQX1 reg_out_cipher_sample_reg_32_ ( .D(reg_out_n245), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[32]) );
  DFFRHQX1 reg_out_cipher_sample_reg_24_ ( .D(reg_out_n253), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[24]) );
  DFFRHQX1 reg_out_cipher_sample_reg_16_ ( .D(reg_out_n261), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[16]) );
  DFFRHQX1 reg_out_cipher_sample_reg_8_ ( .D(reg_out_n269), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[8]) );
  DFFRHQX1 reg_out_cipher_sample_reg_0_ ( .D(reg_out_n277), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[0]) );
  DFFRHQX1 reg_out_cipher_sample_reg_113_ ( .D(reg_out_n164), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[113]) );
  DFFRHQX1 reg_out_cipher_sample_reg_105_ ( .D(reg_out_n172), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[105]) );
  DFFRHQX1 reg_out_cipher_sample_reg_97_ ( .D(reg_out_n180), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[97]) );
  DFFRHQX1 reg_out_cipher_sample_reg_89_ ( .D(reg_out_n188), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[89]) );
  DFFRHQX1 reg_out_cipher_sample_reg_81_ ( .D(reg_out_n196), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[81]) );
  DFFRHQX1 reg_out_cipher_sample_reg_73_ ( .D(reg_out_n204), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[73]) );
  DFFRHQX1 reg_out_cipher_sample_reg_65_ ( .D(reg_out_n212), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[65]) );
  DFFRHQX1 reg_out_cipher_sample_reg_57_ ( .D(reg_out_n220), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[57]) );
  DFFRHQX1 reg_out_cipher_sample_reg_49_ ( .D(reg_out_n228), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[49]) );
  DFFRHQX1 reg_out_cipher_sample_reg_41_ ( .D(reg_out_n236), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[41]) );
  DFFRHQX1 reg_out_cipher_sample_reg_33_ ( .D(reg_out_n244), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[33]) );
  DFFRHQX1 reg_out_cipher_sample_reg_25_ ( .D(reg_out_n252), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[25]) );
  DFFRHQX1 reg_out_cipher_sample_reg_17_ ( .D(reg_out_n260), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[17]) );
  DFFRHQX1 reg_out_cipher_sample_reg_9_ ( .D(reg_out_n268), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[9]) );
  DFFRHQX1 reg_out_cipher_sample_reg_1_ ( .D(reg_out_n276), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[1]) );
  DFFRHQX1 reg_out_cipher_sample_reg_114_ ( .D(reg_out_n163), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[114]) );
  DFFRHQX1 reg_out_cipher_sample_reg_106_ ( .D(reg_out_n171), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[106]) );
  DFFRHQX1 reg_out_cipher_sample_reg_98_ ( .D(reg_out_n179), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[98]) );
  DFFRHQX1 reg_out_cipher_sample_reg_90_ ( .D(reg_out_n187), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[90]) );
  DFFRHQX1 reg_out_cipher_sample_reg_82_ ( .D(reg_out_n195), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[82]) );
  DFFRHQX1 reg_out_cipher_sample_reg_74_ ( .D(reg_out_n203), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[74]) );
  DFFRHQX1 reg_out_cipher_sample_reg_66_ ( .D(reg_out_n211), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[66]) );
  DFFRHQX1 reg_out_cipher_sample_reg_58_ ( .D(reg_out_n219), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[58]) );
  DFFRHQX1 reg_out_cipher_sample_reg_50_ ( .D(reg_out_n227), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[50]) );
  DFFRHQX1 reg_out_cipher_sample_reg_42_ ( .D(reg_out_n235), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[42]) );
  DFFRHQX1 reg_out_cipher_sample_reg_34_ ( .D(reg_out_n243), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[34]) );
  DFFRHQX1 reg_out_cipher_sample_reg_26_ ( .D(reg_out_n251), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[26]) );
  DFFRHQX1 reg_out_cipher_sample_reg_18_ ( .D(reg_out_n259), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[18]) );
  DFFRHQX1 reg_out_cipher_sample_reg_10_ ( .D(reg_out_n267), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[10]) );
  DFFRHQX1 reg_out_cipher_sample_reg_2_ ( .D(reg_out_n275), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[2]) );
  DFFRHQX1 reg_out_cipher_sample_reg_115_ ( .D(reg_out_n162), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[115]) );
  DFFRHQX1 reg_out_cipher_sample_reg_107_ ( .D(reg_out_n170), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[107]) );
  DFFRHQX1 reg_out_cipher_sample_reg_99_ ( .D(reg_out_n178), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[99]) );
  DFFRHQX1 reg_out_cipher_sample_reg_91_ ( .D(reg_out_n186), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[91]) );
  DFFRHQX1 reg_out_cipher_sample_reg_83_ ( .D(reg_out_n194), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[83]) );
  DFFRHQX1 reg_out_cipher_sample_reg_75_ ( .D(reg_out_n202), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[75]) );
  DFFRHQX1 reg_out_cipher_sample_reg_67_ ( .D(reg_out_n210), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[67]) );
  DFFRHQX1 reg_out_cipher_sample_reg_59_ ( .D(reg_out_n218), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[59]) );
  DFFRHQX1 reg_out_cipher_sample_reg_51_ ( .D(reg_out_n226), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[51]) );
  DFFRHQX1 reg_out_cipher_sample_reg_43_ ( .D(reg_out_n234), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[43]) );
  DFFRHQX1 reg_out_cipher_sample_reg_35_ ( .D(reg_out_n242), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[35]) );
  DFFRHQX1 reg_out_cipher_sample_reg_27_ ( .D(reg_out_n250), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[27]) );
  DFFRHQX1 reg_out_cipher_sample_reg_19_ ( .D(reg_out_n258), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[19]) );
  DFFRHQX1 reg_out_cipher_sample_reg_11_ ( .D(reg_out_n266), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[11]) );
  DFFRHQX1 reg_out_cipher_sample_reg_3_ ( .D(reg_out_n274), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[3]) );
  DFFRHQX1 reg_out_cipher_sample_reg_116_ ( .D(reg_out_n161), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[116]) );
  DFFRHQX1 reg_out_cipher_sample_reg_108_ ( .D(reg_out_n169), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[108]) );
  DFFRHQX1 reg_out_cipher_sample_reg_100_ ( .D(reg_out_n177), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[100]) );
  DFFRHQX1 reg_out_cipher_sample_reg_92_ ( .D(reg_out_n185), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[92]) );
  DFFRHQX1 reg_out_cipher_sample_reg_84_ ( .D(reg_out_n193), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[84]) );
  DFFRHQX1 reg_out_cipher_sample_reg_76_ ( .D(reg_out_n201), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[76]) );
  DFFRHQX1 reg_out_cipher_sample_reg_68_ ( .D(reg_out_n209), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[68]) );
  DFFRHQX1 reg_out_cipher_sample_reg_60_ ( .D(reg_out_n217), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[60]) );
  DFFRHQX1 reg_out_cipher_sample_reg_52_ ( .D(reg_out_n225), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[52]) );
  DFFRHQX1 reg_out_cipher_sample_reg_44_ ( .D(reg_out_n233), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[44]) );
  DFFRHQX1 reg_out_cipher_sample_reg_36_ ( .D(reg_out_n241), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[36]) );
  DFFRHQX1 reg_out_cipher_sample_reg_28_ ( .D(reg_out_n249), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[28]) );
  DFFRHQX1 reg_out_cipher_sample_reg_20_ ( .D(reg_out_n257), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[20]) );
  DFFRHQX1 reg_out_cipher_sample_reg_12_ ( .D(reg_out_n265), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[12]) );
  DFFRHQX1 reg_out_cipher_sample_reg_4_ ( .D(reg_out_n273), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[4]) );
  DFFRHQX1 reg_out_cipher_sample_reg_117_ ( .D(reg_out_n160), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[117]) );
  DFFRHQX1 reg_out_cipher_sample_reg_109_ ( .D(reg_out_n168), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[109]) );
  DFFRHQX1 reg_out_cipher_sample_reg_101_ ( .D(reg_out_n176), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[101]) );
  DFFRHQX1 reg_out_cipher_sample_reg_93_ ( .D(reg_out_n184), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[93]) );
  DFFRHQX1 reg_out_cipher_sample_reg_85_ ( .D(reg_out_n192), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[85]) );
  DFFRHQX1 reg_out_cipher_sample_reg_77_ ( .D(reg_out_n200), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[77]) );
  DFFRHQX1 reg_out_cipher_sample_reg_69_ ( .D(reg_out_n208), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[69]) );
  DFFRHQX1 reg_out_cipher_sample_reg_61_ ( .D(reg_out_n216), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[61]) );
  DFFRHQX1 reg_out_cipher_sample_reg_53_ ( .D(reg_out_n224), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[53]) );
  DFFRHQX1 reg_out_cipher_sample_reg_45_ ( .D(reg_out_n232), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[45]) );
  DFFRHQX1 reg_out_cipher_sample_reg_37_ ( .D(reg_out_n240), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[37]) );
  DFFRHQX1 reg_out_cipher_sample_reg_29_ ( .D(reg_out_n248), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[29]) );
  DFFRHQX1 reg_out_cipher_sample_reg_21_ ( .D(reg_out_n256), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[21]) );
  DFFRHQX1 reg_out_cipher_sample_reg_13_ ( .D(reg_out_n264), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[13]) );
  DFFRHQX1 reg_out_cipher_sample_reg_5_ ( .D(reg_out_n272), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[5]) );
  DFFRHQX1 reg_out_cipher_sample_reg_118_ ( .D(reg_out_n159), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[118]) );
  DFFRHQX1 reg_out_cipher_sample_reg_110_ ( .D(reg_out_n167), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[110]) );
  DFFRHQX1 reg_out_cipher_sample_reg_102_ ( .D(reg_out_n175), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[102]) );
  DFFRHQX1 reg_out_cipher_sample_reg_94_ ( .D(reg_out_n183), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[94]) );
  DFFRHQX1 reg_out_cipher_sample_reg_86_ ( .D(reg_out_n191), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[86]) );
  DFFRHQX1 reg_out_cipher_sample_reg_78_ ( .D(reg_out_n199), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[78]) );
  DFFRHQX1 reg_out_cipher_sample_reg_70_ ( .D(reg_out_n207), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[70]) );
  DFFRHQX1 reg_out_cipher_sample_reg_62_ ( .D(reg_out_n215), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[62]) );
  DFFRHQX1 reg_out_cipher_sample_reg_54_ ( .D(reg_out_n223), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[54]) );
  DFFRHQX1 reg_out_cipher_sample_reg_46_ ( .D(reg_out_n231), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[46]) );
  DFFRHQX1 reg_out_cipher_sample_reg_38_ ( .D(reg_out_n239), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[38]) );
  DFFRHQX1 reg_out_cipher_sample_reg_30_ ( .D(reg_out_n247), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[30]) );
  DFFRHQX1 reg_out_cipher_sample_reg_22_ ( .D(reg_out_n255), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[22]) );
  DFFRHQX1 reg_out_cipher_sample_reg_14_ ( .D(reg_out_n263), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[14]) );
  DFFRHQX1 reg_out_cipher_sample_reg_6_ ( .D(reg_out_n271), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[6]) );
  DFFRHQX1 reg_out_cipher_sample_reg_111_ ( .D(reg_out_n166), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[111]) );
  DFFRHQX1 reg_out_cipher_sample_reg_103_ ( .D(reg_out_n174), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[103]) );
  DFFRHQX1 reg_out_cipher_sample_reg_95_ ( .D(reg_out_n182), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[95]) );
  DFFRHQX1 reg_out_cipher_sample_reg_87_ ( .D(reg_out_n190), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[87]) );
  DFFRHQX1 reg_out_cipher_sample_reg_79_ ( .D(reg_out_n198), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[79]) );
  DFFRHQX1 reg_out_cipher_sample_reg_71_ ( .D(reg_out_n206), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[71]) );
  DFFRHQX1 reg_out_cipher_sample_reg_63_ ( .D(reg_out_n214), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[63]) );
  DFFRHQX1 reg_out_cipher_sample_reg_55_ ( .D(reg_out_n222), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[55]) );
  DFFRHQX1 reg_out_cipher_sample_reg_47_ ( .D(reg_out_n230), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[47]) );
  DFFRHQX1 reg_out_cipher_sample_reg_39_ ( .D(reg_out_n238), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[39]) );
  DFFRHQX1 reg_out_cipher_sample_reg_31_ ( .D(reg_out_n246), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[31]) );
  DFFRHQX1 reg_out_cipher_sample_reg_23_ ( .D(reg_out_n254), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[23]) );
  DFFRHQX1 reg_out_cipher_sample_reg_15_ ( .D(reg_out_n262), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[15]) );
  DFFRHQX1 reg_out_cipher_sample_reg_7_ ( .D(reg_out_n270), .CK(clk_48Mhz), 
        .RN(reset_n), .Q(reg_out_cipher_sample[7]) );
endmodule
